`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
KmaUx9VPc30mrkuCdvJ+AP4qrQDYygs3MJhQrNtirMQVfAaZqCRk4o7fVqXkEkCp26yvFwiujzc7
0V5BMQmfTw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Jih+r4fiEHZNWQYM9OpTmjyAMKKS88l+lni2YfMWRAuE6jNNoDVkQyMa0CWEBiqDlUdb1gJyphVI
jVncJdi+3PIHXTM6c+tEehu+eVV6FvBvFs5BNcmpuTs8hOzN/4YvkNLFd8fWWSGuQUfk9h9qu5xE
lakPfD33j9DKd28JAl8=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
LNLNze71NwclsX1An4C1xclzykLXvlLHF+MaaTXYFQpTUw9M8FJZPpPihy99JJ5xkIp7crXeuf2z
XrlX7zR7UKq+R5jc3iNyv2SB81M1SBWpfsrAvMtVwblIa/P6cM/i8waLPVqFmRJ/UaRb532C4gX1
EyHsW9tpPf8WDZE8bOw=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GpazcOoT/5ZNrkwSybcERaKokkjkNu2noEMgOzB95yiQUyg27+n2cmrCCC3RTqPc5wc3GXo/xtX/
E3C5Egw84ynR5IFplelVtNR9ZDc6bELtpFBurii0wmyBxMqoPX1jpmT5DJNIgjdZoOIpFkiweqUP
iPV0KJVD8aL4ph85rbWIU9YTHa18s2h/1dVSmxbYLh9kooTXgdDLOnZqLYRoXuBwnZ8V42ItpAgL
sQr7yY5JorXlsIHx6LmoNXAGcdujt759NTVi+yvzB5qAY8EvV5zCKu7jBs4It6WqA4fQd2BaqpfL
wj4QMJpAPnkceGNyhfLsU+vIQ8qzLhNq4iLl3Q==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
XkeXYDKAjDl1eSJrgFaRJg2i9bWQ+LkePYLnLDHXrmf37dfnoYNNRhPB7rRcZXkguVZwyvmOz/1L
cQ/0FsFt5XiV7Mrse27uMcjPCZikdAAmqZrRCW1qCf4WuDsw5Z1tCeysN0sFewLQ5edp5bHFgLyy
VsY++uVhlymgFMaiLeh6QLGh+om5z6/2RbZBl01qh17fBvTaCkl8wg/YiBZfvY4emkxNVevGOtjx
BJi0++gEMOwnJFnhY4lens/Qp+LSieFkosckHt1ycFPHzNTz1Js5sfBTksBD0IhpHnRNBem8bHZb
AM1YUSCwvat+ga9g6XO6oZENj0bdyg9fKGqkzg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
V/rZ/9RAvX2gj5U00mVm3EF8bRlWglBkKdPzUohhvVB2DZJ8WEyCATElI0oAFWoUkJMHcBsN/R3G
RQtAlO+WBTAKpNrAhZEcy6JLV9+UbOMb2ntzKo6hmwHFdU5/gYB/f1FHVsWKTk9edmMGHFEYJ7Z8
4x/oPFKtAEnuDJgiLSOy6cODcYjhsScFxSD3Il+cLvRvwDfrskzx7n2d4h1OHWtX4Ruc2ijj7GMT
aqNxvlQKqLaMiPnHjs5+orSA7aREva64SwnXTuZvyUFocsQZnZqs4rSC0Z5rXxRBdjZCkN7LZEQz
Hnz7H2ykrV7m7K4DqjLXLKAU5Ea2P8R2NiB5zg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22944)
`protect data_block
u2mAGog/yC/bJ5ebYqeFyux5uuufhfSHOr4k6iVBsmyW5di58yaIE+rHf/OVS9aVjW6BEj6DY+th
sxkb6y7cBLZAxIwupimlhL7RpJAPS7lV89J/RIIQX6iniDiBTBcnZoutfvOL1Iu56eBKpQVVUyNA
W6PT0ofgi4CGDTCE4/Li/Omro8L3rEpbZIsLghtIj9jzQgorEyvDOralLuiSXtAjPtLHUSzw66uc
06Mk5lyLlHqPa7N6p3I0lvkL7QhR31z60xhaD0YOfETIvILKU9rxKlxEiKTlLBjeIvkdfAXPQd0m
8BzsKQzx6CXuyPkrHpLI5RiRMWOm8i0YMuRTGEuqYOG/JbN1q6xpeQz03u5ceL/zkA9uHiVMbbwM
xUDGiJoBD4UhJ5fhYhA9QL6EJ3DeAfifc80N7ZqCtg6BFPWQvzU2ME4M+Ep0L1YIGJI4sAQeJYP+
+CGkdTuz8DY2SzjHyGZ6ftCjQkt3pT+k5rzsfxhWrF3pFGI5lMZTsBYE4kSKOVxNenabnYzJIMLC
CYaEGWCxsGgLzXPgr31S8vRtV/KjTpJsUqfEyWVAy1WlFMBdhPrLpSO2sWJpwgIcdTCfZXo2BUv5
4DT0KK2focxAYTWWqdOnF+nk+X0o96ucjR1Y5PMOSbMjBg3hsjIKuX8GAt41LULYWP6fUHq7xqBk
Rke9N+pBkcaULrVE2RwcKYYh/qnEL0kj/AEUyRxKP0iQc8mlxNK8gElivAsJJABM4l0FGRVBkDO4
LRKbAT2ARStyMHr1LbGZ7vxFAGupACb+2smyS7oPZ99eXY1Oon585cppS6Hj15icDXETulNLR8WG
tQzBxYyWBYEImKXCi2ZcCgdLOc56Wk7v5uGBdvbaamlgD0lGOEFHD9EprcDvi3LqBpa8e9V2U6MU
zPV7zyC4RWNdWQAPx6rGTckm2LIQUI/tFilzdIJlWNXFlMFnj/RZQANEULOqggrJSVqd8mUXsAIR
G2arp/uaegrToBC3RTnkn4R8FZU2Ta9Xn9jVWeawE2xiPnUuoJbgbvMap7HLL4/T58nahC8mH/h2
c+4jJrSdcsnzdzzH2v2W4FA4aZjelXbl44ZCjKyErtP6Z8fq1cM5Dv8WV/KplSZxJdKmjeXoj+6V
kz8+OXwYruMWubIPtUOcnyW5N2r4YrfQdnRNac573PCUm1jVURg58pJyrz/94i9GbWU5BHCjlm2D
ym5OBmNRqkdvm7wxiEpz07504Fo1DxNP3PfWISfoTiPE9BSo+1p/qZiqk+CDs1Um8L9nAs+wxAdI
GnY31RIJUaPHm7T3cR5F0PnQAJ6vRGlaXk3Q9L1AQN8gZ69BJysHuXTePPPWhWh2JY8g+/ATkPkO
HPjMTTWHJGWOlOObhM7LWLYtTgiItI+74cxBhbQHufHTMJjyxRORvJ1w9xNUEBkcIDrdSUTyb4IV
KdAZ9yv627EmkvoHtxrGNFcW5ZoT5IF8yx8GaGJ05qR4FRmZjKQT8cPLyLUEo+8+LD+wd3/5akkS
v8PJXq8/o0X+NtomoWM8mvr1zdG3/x6ZhE09tDJUPgwdcjRnjbYk5GcG8p6dJS5ZiQXZSYdORQja
GRf35LOeLJNFbJkyIIPOolsVZkabbv7ZHayomNb5ujnqwu7zAtd7Fk3cSSQTqPipULxy9tdoku0A
KRzN1L466q2PuFjHWt8dX4BZsXBdoIB+NHGMIvTxEm9Lye8/AfnZajCj1DaxhP1IMU+AOZtwi1+S
qpmN72KwagC9x3h4vlU5yGHEkFhQ8ZL7yGzjwWS8c5u/g0kIz0EUJIYDPKB0sLbU4iYH7jbOgip9
krcJJs67yYwJh0U9MLtE3XBHsV4xPaFJ3U9hiKl1oMilIRjw+vjiR7bGeJ33sNxp7Kn81K8T4JRn
oRqm+VlOHQuQNAV0xmjxBAyo42RpXaqxRKZK4S3lP4dKkIaSkLY49jq9mdG1lVsFoG8fonl+aGyl
8/RUfPQWSmz8Tt8QOICOPJQLkvjmvYEYRPa6az1QsDYCgxPTY2LKYcds28w3H7YPov7ZO4QgGc0C
Vk+HZBLORd6xRyjSXmeewnqfDJJQTiqorzA9RFYvLFZ60rMZ8UHYExqLU8q8eN3Xxs/JtMbjqTGL
DSoqysDgJUWoG6gWQGQDyiNxQKuGOCzzOnAXh+9b1TFl+D+/vQfgqQSid5eZw8S8kGW2zutb6t4s
tmegrOzhVDVAdix6PkhOgFByGpj3anyR7IRHdc4aNH3NxHNJplRfL2kCCkJIQ9qeKot9QmOoSQ9S
pfm0pZEqx4te6RIGjArJcx/+b1+kfYh0e0lY4hFvzwK0OCdOVJDpqxtlI3z/mPg8A+IseI0rAUE7
D+mb6IP8OxkBhWYDc2sllIMukp06nuS2OsGa7K2TsFZ+7K0SjWSKXMCsQix4LYbdYC6XhF3i4jqR
XpWmLfPwxrg0YyvQ2yQPESlA2Yr0QUOD2aHBQzkWs9L8WmlnhvXIHOOKUV+IVoEpl4uLdbMu4bYo
mgcN28ZiUu5A+9g7vDUHxa5onMGlpRm27SHNbQ+v7RJHWLkvgPnHLKVZ+x8PdHK7seeGiCrc9zog
IsNJ3qp3/AxnbYjt/Sa5VUPiPgg9g9qV96g6jQB4aWAJS3rA0yP9nkUsKCFejmveNSptJrDLCzem
3I2YnArdImJJzzfUmc8K6P/5RN4FODuj9STz75sJh9tCaLP5AtGHkrKXOhSEvmbqrL9oN9mnEbZQ
KvtcNXDPkTUzFmLJkHtWdJTvZXVNz6fiOISc+GAPedNLf0ABKmofa0bAFAAhvF04wNXXhcMSwsxf
8rdgy957mpK6iBFOSz8dZPiwLuf7/Eq1u096CphBK2Zm5vJLltekfuCC/4aRXxCSUgSQJ68tnWAY
mT2/hzXLd1phAfj68j/wtwgdJVDt+WRSCz0BMtCaBq/If2cwgwfVE2wwbQL5mRk5O6p05dad1CBq
xtD2mFRzv0qh2Om2JZPsqlBjLbjbi5OfgWJp0LiBfRtExRQR8iawOiKm1QAPORENcyxMjDJIU4UA
LUA9fpE1knym18AcRZ/+u55R85e51aXvUr5vFrGDB69OemzVBz54dU3JcYhJdLoZjGvCJcTYMYgY
IZl9f4eOFK2lWeS+Mld5uAgYFtRD2HkGqOZe6muHGtCCVY4qBC4QmU8CVG/LFPLcaRP4pAmpWBOh
a5PcgUlVqjREfasEHQlnMFKiFUuIt7P8Tgl0bjJIJcxaJNUPpxmodyeT+uijrwqRb+6nabjdwVoH
s2X1il7TEDyYU1pbqshAESaUc5TGUc769To9WX9MuDfjBwSJq4CYKIieA2gy085PG7SLAswM/oif
xV9MZyw/i9wpNEsO4DUC6haGKRXq14kckwb+0eq7SBpmvNPxL/NI+RDkzRhBbG2R059ELpZQ+Xc4
UccBp0T3MyzbLRnpEF/IohdyJXbfnoctb4UVk9qQk0pYfnsNWdgcbMQdhhruE3L6kiOjj2eaXap0
bUMSIeL57ila48km8/B7qre7eacw7y002zMDWnG0doIfc551J/r3MXttQHw3XYBARt9RU1zUHy6a
DEiiGzTcXMecLvFNqLqdFQVRUJaK7rPIaNMaEHxtQHogNOjHXNhx0GCNkVUCkDPlRvtM6Ca+eh9d
xqPUSavfXV3fTi3WVYpECJlPgHJ4lGWZ/yVkT+H3FdphOXAastQ+fqGbR5jOg521ziQdZL9254/f
zoIzyLRwN807atqki+g+k9sOpwxXVc8mP4lKw/cfupGI6ZMTXWsvri4yAA4koA7ZmFjNdKkiW0/0
24C0bs1y/r8WovAWreRXRI+e1Q0HS0fTgIHrL8alz+gRd46Zkr3IJjNML4Zr+vjshd/Wl2ubXFGY
4a8wdKKc780AkdXeryNa7CjIKFC0Nd1cQt2cHZ4sFssTjzJjDxM0M2Zy72b698YSxvQjI8IyEZxn
epX1xvbX3hBPVboAulbjcbtJfVJN8BOpZ5BCVo7NR9lRdbEszlMrrq3BME9iwMmAbzkda+y0rP8I
KBjwFUf/xVTBQrG7KJbJyBFEs6QZLSVCOJZyDd5le7ZGmYA82aPknUi6X4gm6O8u0jOBhafDoBMT
qZvLmoSP00MF1Jh979gv8PQfPNyMPIPnyqbEjIFAydXn7gteCsU5Z9TZHTLiLRpyJ4HxvvNil5FC
L7tdHfubAn0FSyXDaYHbK8nNjj6+KZpPQpum5OM0yK4gAq5aSKzGq6NWYJ+JLkadOZx44gWhVwrn
z7X97GL2ZGrf+pVSCEbmhwhuB0AoFeY8h7CIpbQUP4jXgwGpLK5mOb8Kex3nUsid55WmEcYc3/IE
SLU+ZjKsoOMsCk4eIF+k1+I+f4v8gALmwpadv4Y0S2ff8NuRPxVhG6MyEXbZVBrnX0tRlHigoAbv
3JvrUjOADu5iq9zJsKvis1WPCg5A9IcwT75GEJ1nXRrxJXhr/0eRZgK0rHbWK4re30ZD3EPlrZZi
iIBAd4f0g4zw6kdyR86l6Crv5vCC4o03akSx/ZnUrgZa+UBtouNviMgHCCTnYf+1XBePb9p3HJoj
Y262YpUo1dxx9a+EFKE9vRbEfnFa6q5NSxmHKhKppS0gdC2AcX/jjVz+dyua3d8qqbJG+x9XEJCx
tjY7kXVDmmXpicNYAMni7EltZZJ5B4nuEtAB4kU7vusOWboj891p+YGi7qcr5OtstXFD78PzVEf5
2qHgCU7vJ+AK/9R96hF55wZz/UdJHajRYE6mmIlyBZNmvJ10c82QTWg6SXAOmfKnCurYTYII1/Lx
D+jhJ7SHG7SOTa1pzQIJLnerFVr/FAPX/9alr6J8HXbfJpUIYNI7MrVQdUeEzHqWJBwgShRNmzGS
BXkEXzDQVHV9sUFwqrS1jv1LbpLxu6xrtyiV5x2UFauTaaenZOTeQnVSoVRLTgEu20ZFn9YUcSIc
pfFh5jIFiuUiNjTwR/K0FE3MS2loMRfuttnmmt+o7VWTb2Q2SkLCv0FYNFwW8ZCK+EUNTHKcg1NZ
9UafE/1mIDwatq5ys0lX9Dv27eklx0CXNlovrc8CbJL9Y3scgBm68TPAj/Pk3U/X3xzpfwSrpQm5
KSyM/ATKckOOKfW3/6yinMp1ShboOWw8GYvtNY1Upgkujzrx1pyZ4ZJKBQo0eb/CGwePkGOzXLze
afjSOJLf5A7sixNVzQ0MML4Bfre+pmf75xraAz4f9nXM3jC9ukk12pez2Ec3sqddT2uwfUdBiLfl
hoQQ3Ic0nfMLaYadE6fwpkBWStQd+lVH1dVtxcjIqNJTf6VAtpLA35aQV8hArbtmCscCc7I9BORK
6srADiv70Eot4PGk3GnfutMBtiOv13N+KBO6IZEqC8whGF5+Lro1nnfk9m5UensB76W9MleGYeHj
b2Kk7x0zGWpS1EEGUl9DqTTxnqUrhj2o3q28b/BcGa/irH5o7ybLPJEPdYe/XMKtqfPYziHEgSB2
1T6+6TOqOYWtQtB+8MVXUxEiD9zPDDt7n07uot2seAeGXe/WOLqmxwk4osTUL/3P9JDcV2//m7+i
OiX87gFNnJlxMPkLOJ4StWNfRuWKokGJgT/CR8s6mNufTJ1qpwNAhNb9D3mwmAAw8hl2bsT1Qcp/
9jmTdLqwulLSFF3vcDmOWsi9ZCy7IqLDC8VNf7/flOottLN6aFkrvHKwfl7g8i1de8DfaYosDnAR
3v09//HM2fLsyAXvGnApj8529FagIuu8SGZ9pyGspFDSUPSQqkBNxjKVDsmXAshs/+ZASaxkmxOz
tQRrgxMrbfrmoUrOC+GbrkS3HHt48eiqC+OJCeQ2v24NDVQGgEbPrD8rpMGNGs+xP70qThiRI/D+
fq9PjUt7n9wyRpd/rPY7KQINHlhZxeWUHuDSCDQZftBh65sERvZLdoTCohZyalE6AhT4Yj7GULiu
AOh0oglmjWHMynTP/T1w9ppBABNcPsyYnlcnR8OxLD4+/REZS12uu9lAGTPgphumktNNSu9NGocy
eVpQSRt+6q5QQ894D/Tedlv505g7flVoNf/ynrebYOgEpnTL65k8zUWvsV3KlQ6XeHw4kcdjqv1E
rVzMii538h2XTGNQa+n1i0mlQkmeiCf5UijVucVKOtEkidmdZ17qLdJD/DbSR+KEYjXMkdP9VVJJ
LAxFCDdkj7eJRvdiBLT00gWYOEBLYXlf4uNFYOysBnEYPS66oUUxYyKFm46SWDySlNDyWxm/zcqw
NkSUJVBcshdi4BrQXRJRk6HP88uQqqDqfqF4VV8gXnnh0wBe/hcRPQGshkphffUM9zQlevff29u5
v8jgjmk2gY35GNshLFBBKEIDY/tWAggifnEtieP3BV392ZNmfSkwH6fAAkvV2pC+bqrMCvB+hiCd
f1NOIuosMy7WKX7A6xHMs+s+05dhdHZYU5B61lHWJ7qagg5ENt7LCFY9Mi0nSGregO3c/+NCwJY9
fCbwMfqa8hOjEZvwKtMO37+STERWr/WXnrS6/mwj9UIjaVzBbJWed9bt/YYARN3nB5GJvTG7Ad4L
gVVCVBf1cyIgiPcvtIfYsmhSheTJfG+pz5Nnz26y+U67iLpU2sSuD7CML8tijeTXTDQx0zH1H6j1
GxrXpa+0L2iFWRP0TKSqkigkj0V4UbV6cnF862lthNUaONSaOzFhZ9/XxpNS/9K/AU5Jolw+D+9R
cjWZwbKOUoxNvCY8nQx3W11Tgf1egr9C0Oq0wb6Et+EM4ZnVZlsWvAouct45JKoneZJP/MKsZZUV
4SSojgiLP4Ehea43QZFoy1B2hG9VniQZsly6YrNcRjS9G7X+MuzaeWfP3w7BzYUnOSewt/70twdG
yQc93upPhQhwtYBWxPWJcANqwBscXOzNVG+393bJzCDMBwbIWP56ykrqEFPUL5zXo8YGNLh6/ZxJ
zZNhyd2qm57h9HjKnN5fCYqNB7kNhdYKEAhq9FUSM8/WPOfVPEYLxqoBkjMVexIW7T4yobCpyU/X
OULlRImJjxvyNSYXYdGRGkQ+iIro17Vavaw+hykBWhc/JRh0DPUpdNzAg++i8qR6FeikbyIQJ2x4
kgYzIFCE/+E+0Pcy3lAXKaANI14095ztXZBtu6ejZ79OebtsSgp5yGudXoW5c8f2VXGRU8CoWaNe
pXfN051POPsAK9y7Hg5nUzoWa45qEIBN9u0GL7dsXNmS/5rQuWB5NthUmDRcXH6zo5c4XpWEBWss
7VlOrrEysdunnHtYGJFnWbKQidWFhrLgdqz3VLt/HAgEee5p95ArUaZkK4+xadk8TorRlNaTndtr
9dJQCCih7puOUO7MJWBfKsRBsIRPI3lE0+mMMk5t8VtCAYu9EsWPq8BiQGsr7tT5i2775JHLYFv8
U6kOThwNUzkILFguxe6dywGAd2zpZloPEW0/TG/dmpCJPsI23rKs0sSCUmhBiWz1YhSJHQUAl/Z/
kOuth8ZTlxntIMr6zLcbsML28uwVnfGsGShU9Y5H9+LVhrEYDhiMcn0/qWhnCuFwzZDlB+edNLdK
gMz3s9JaEOpAtAk2RvT74no2SjB0eHPJAqjgsinuDNHI1w7poRefbH+oADS09gACmipmZKFaQSuv
6Q6qmdSEkhFgaY6S4aLsu/to8QE6b4vEIQnk9rn01PBMSNwGwzjPIwKnpKLelaFHs4sOLzOrDdU4
veFjURVKcKG3Nb4QEwwU0fBOK0mxDJ1ZIO5BpDqOjNh0Gj/SIfOfbVSPug6A3e6lank6uGZEHloK
Er1AJDfPdDu/UldzPJr484nRJpjXp/thd+HZyhoMHiB53Rz/HK7xJKP3/L5zEdv5IdEyRKSyaXW6
/HfAaGV6OrO0G5ynDCIAu10+USXTP/y7zMt4b6prGznGDws6y8S4/hQVuLLOJZtuHqk+10ewcyx+
tG+KO0ay4tlksr/Eea5ymBGoNUbaaezBNJkXkUjU5zVACxJ5OtggS4SmrQxrLfbbY3QxdoHqMSd2
8S/BuwTzw0vS4NKlx4bcT0gpl/GfvURebEDnmjo19yZTGk6xAx92gpNI/OEm9jEeUBrUHlO1Hxje
Q2YBOMIdmy0EZ7Z9qiwiaEltWSYwBtj3YUoFUR2KcF3CdO9LV8YPs8K/GW+W0Dqtf1slYcl/ozYN
QXLj2NczaCy6Hq7YJLCK354fH8/ZARTKGnjxiinWPS53++lZpR74zV6mkb2hysoR6sSAB68nN7An
t5d7YgWViCyVswJDcCK2U51uyZ8knPSTGuWJdhNyCDCNpW/tuEp7KXWD4D7JeEoQ6oRsvYLErZI2
fgRnJONuwEZFBxxLwFRVnltzb3j4TuGwr+T2GfNnJ+3ctbqK4wn2qpze4I9Uz8tNBK/ufZ4TbQFr
F19EFFv2smKVaEqUhxdQWt4yxffz9LOtlRjdEiDxAoHYdXeAZpKQpVXY65C9qXra9PUNThF9c8e2
oniDeqDkWT6evHbhdLV1FiErJn1S4Ocba61sNa84+3KPvkd3w9YI2RYIAnMQTAwBLuU5EW0Ajlde
LQV2dfztQGS57PXNRofEggHWrqix63k0q+NpTu3lPJqKx19xXIsfXt4OtYGpluEVOCtI4UD++vpD
C1zIUuZVD9znoffJ1NEjvzEQ0kP9z4uoCFaWjSPjsQjnX3Z9RaSq3E3VYEbWiuBIxhh+wAIksyB/
rA6OhQMRLMi3K2a51hYjkIsBqzfD+Cv0UQY3+fDIjBCUsR2lcJRlkdyj9PzV3kK34yemiiNGUrCO
uOIHATW+DLNrf+rjciuqMqZf6DzCgAy2NsopGlBg0mFDSDFW4s4MaskwkrmnpkD33Rx8GEL8yQa5
lcSDldKmqApMvGbtJah3vblrSFBf/pq7Zga3w0urf8kJ8qEOPGvNMTnXA5nv57H8f7gN323gbADe
Aw2elsmhcIXI1ok5tnf2+FPnJAtW9+119IOMKewLEO/MPPpdORBT07D4rsrrKvIkeSfORZVptt36
Bjo/gN6y4Ppdo4wB/Eu4lQem+0KZ+gaaGVvoa7FYIR+xUFUw8NjFQ9AD7/2NNZuJL9J+IWE8quP+
NW3yyJvM1mVa85tx3bJYf5D7fY6Ud2wzBNWQfprEafsrzvAKRSZ1bnu4ozeXUgY4EBx3RPl/D3G5
Y8stEkJqT4pLrXn442SQWW8eK0o2o4tnw4fYZLLIOUQ4WYbglnc4ibQwGBvLcYVJn8pk2fKoxUEP
TNdsMrGvf8aYgxpC7M4F1ohoix9n+wWu7GKBaznU7tWze9XAonBGId29zcCpZDf2KY3cahBru3WL
ibW0NAGQFdu5qVM44D6Lqar/RuZ8j70HuvYLsfBUR6O/NFgX0DshnYLRA3vgxVPNgVa2hLeML69p
htfuZV5nsUAqWmnsB9p37mybvP8Oq01SNJT/xAJA7ak/mKsjvnJ2uae5lG1Hvk1DNHmIifAAxJtS
hvIq27QC6BG2wtFIt9FBsimwg5WnUfSthfFp2zXzuacky332dCcQA+aBOT9qR9ZI5xwyUTAAlkKQ
Ym/Z8EH1zuxTkAuT33b3cHJ++rej2oiVAnG4DrlCKwD0AdxAmBqpgbDaXeyPOkqdF8syqPuuAZjq
Rxuq7kKr/5lVx2UhE8gZstXTCj3QbavCLc8RrVV6WlfJzf7/jifj8q3YSQVe83e44L7osCCMGj8T
Rm2JljQITTgSv4DnSOsBpGcNGS6QbzMNqrWqGNYd7K5W9PeLlHsC9xu9e+O8E8MxgTpBsp3+xrJ+
YdBTvAk6vIEv9yTMSDw56UmZ7fNAnEUSGfWg+vBIHR8LKBFvAA7RroOefYL+Wmz7/LNA/484N9JB
01Bt2u6mw037JUs983xbTjcIe19tnIJG/Xryu98GIZhgddqmA1PZijVRM1GyLAICrs7nn0HChWjo
3qSLKqRuqhgH67Y/cmk3z4RCgzZXLkopEopTFQa84+ffDaples6nany8Pa8buOlPh7rllB8hGiW6
BGCFEJiRm/69oDIS917/2QzDB/+xKXgP2HpfsoFFqfjr7x27c0sv9Nruk/y30XGA8+9a/8Z9U0k3
FxuuyN1dr44MY0zPWpkNEXjMbzP7vbsveah6Gab8ysF4aqvk2/q8+2ignbIpJycjENx7S3EFmBjY
/R/lggqqKgswv4tde2KcjN6Zf6UMohwh/xRtg1laPXqhryI6uXdHDEcQjnyuCh90GAuuj5L70Klv
WafLv5rv24RaBcfEzBjURhr6SPS7PH0Uns35S9gDFSHua3xWDp2n4GZ9bJqaimnBRcDUF6l4m/So
oOzP5cUfUtWTAopQdqP8HcSU3r+EfZYJch39Gfda4+r3R6rxbDTij94TyXnAGqhE2IgcreDFFBxU
NlQ66fKrjW1DQ39dyXFJrP9LOUOorM2K89nHnAMcOfZgAiFM+kD3hnKU0970El1tUNLGhhdkJ39h
keod9k9/qQ4+Ff5giT+vDlWofsXRP6rU7gWu9Nbjof4L4U+GWxUd0VySBKEjW7fk70ShxL9PdyXQ
VIndC56As7Ag0MeaWomo/BzKSVpZfIU7a/JS2aB8lIoiOYh71wTwmNoze7n4A7We154yH8WY9buN
QnL0+r/65d8aAFikEJd+oOotthk4TfhLzRHxlU9NeAsY7aoAVxHMzBP3feQTtRQdEaOPXiEHE7a1
hCgOMCQKW6YH1NnLE3DzvDA/DfO525G8Ft9JDUcaHl9bfr6oSkUVp4LMZ4CEHQymT7XjcJvYOI1v
HKVFtUEpvdTiHy+IWOCX72lQQ+uuMiEt7I1gWctY+61RdvK2dnjjEvFVLtMJUaaD0nji+AayNYnl
TNmandq5SN+T4briEWVV4fi+YoFMCWv+Q1rlR3fu2AmQEtGsISrG9y106qjcx2j84U0eeNJVnDEs
+bSaRoCDvwLQ1Y1wbdiCbUo3yqcC/b5ehztXAmWVTea7SxINd6OLV/ZZ9Qmqi2hMypfkPXLAO+Js
uSBJP4prBZi4T4vBnma7g7687WVssUkZkAz2Il+UWfDam0CMVoW2fuCMRyakBbCmO4acFq1tVaxR
rGfapJ7ED5bgU2x0Rn8jz1Z0MT7QtuXpfFryvSWGTI0Mtt8Ms7zwDGX1OaHDTnlNLKpttHml17pN
47VFAtA/+LLBglSi1pVZx19EcoMe3xVPZiO/NmI0FMwcc2N3UbyM3bXw75QH/INIcyvJ2qtiTsEf
2GC2Nt0fgH8+qKn2VZUY57JuxyJ7KUpEknh6CwTKZ/4WaEcUnzoehYWClLVMc1YmiqhQ5/XgeZqD
DRJOFSxzaNlWGZgbkOu6udgSDgJ+d+GjgFkB7u28Ntsph311ux7ipNvbDnI7FFsxe0mWlpInXLqL
Ux9YSxq88mM9ZGTjcKDYbs7tVgs34d3XZlz1PrUefjdOhu5ncCdekvQdB209UhWdO0ecXOUNiOMq
Bmdn8sN8hPulNJPrQcVa2SEcTL8osI9HHFkx+GgsK4idv39QS1ehCoGVgCB8CNomkW680NU758N7
mVUxfNaeyvdKgQvQSUbUfvef5A+mUCsUdei9ogytY5IBvXqLODdTjseIC20c7HXD1inyXPLl0a3u
fdZNtUaUSXsSFepYMASm4xNh7voYoi4S5Omb1gpbTDEjgmE8FTPGfjIso7gCvgw7iTFg8T0SJ88z
/oNqGUKWo9VSxj6Y6jCBhCyQkpRmMxT+SYH77wFMEYTQ/fHCoVqnimdsyWbOWfmy/9e4XR5EtM6L
xX0UhzRXvmJm5NIcrx0qkQhECe/jnK2iNWkLO7Dx9uADAu1U8+S/1OX1JJ9EcCzrLunk73lTp7aP
nr5sH3NZkCkWrTRIbxOrtM+H3XqEMYzNnezLO1Hl4XLL/rHy9rKeFh/V8Kxwhb4MDUoN2cuziSXk
AB+F+StEUejdOg2FRaIUQJe+sCwgxmTUVzJf7qQ52RY8E5nJcqijWS7p32uaeW3e8ZpFgPosB6tW
HSymDcXc7NC0G2yGe6h2SEUCuh+aZ0B24nKtl6kuUN7RS38CKbJH37yloGeyhXvOUmys0EhEZMbT
VVab4/jx0F6Egh3Fl464nI4f/uUrqo6oI8zTkToJ9ByWjrskyzM2EBdgcmihULMeXTRMnZ+smhE7
P7WmZshou/XIAP3w2cz3B6j0x7B3SWfyB1LJ9mBtVnbizD/uluWmsxTZPc80rv6cJxdjqczG+QIl
r+ORKs0jT8sFBdD1RiqRZOCUGQeHvCjlhCoPZ9K9L+DOtWfwhLYMK/4kcKjVCOIKmt/mo+/EwlUL
Yw3337+w+lQqRnmMoLv/Q0DTBVaDnJmGG2NSkNq53lONcnpg+PFqLOQGVeivqgI6VE3gIHCSqF08
og2047uUnR+YpjYexSQiwEYREuvcOILEOyZPxb9kNOmEBQxDF8FwhZel8LGZ7HjdBGC9pMRV0agr
5b/jCM9lG0Ms3iFsfhLNKBS2UAa/xb7U6i0MecilIYRG2EhjBcIHq8w/CpJcJdWIvwh7xSRsIGyL
O4kbIdVRcRIbjyPER0/eobCQEKZwn1WFQVRZKfw7j1L7Vuvj6gAKxoaORsJR0qy2kLrf5mKXoN5e
Bou4WILhyA+5gm5EYXvDyJy5dJ/uxQAUVRC9Lq1pb5M82LbSrlk26oRSQEzkiS9XVLjBVHXnTDeJ
XzUmvz3BQ1fOP6X/AmV9dFd1nX7QTx7eIo2aIwiQ1eDDS8zs+XIGfgMZ48/fElh8lsCxqHSXSCqs
VGBqfx3TcQDN8jW+RY2McgZ7Lu0uq6/r0DhOp/QwngWKvaf+Tjr+g70nTq5HXVVyZ70j/DmaKWu+
+vtghCnLI5h8KwlT7Cyv0fh+0J0f2CPJtMXttsnlzdIi+Iw0ICsMco4Ke0l3k3tri+akAFvkMjfr
y4HvvjbRYsLzd54yK0A5rsYfJ2P9Z35sqAOc4nrkSGMGpz7rraU5hqdt/SQLrs6RDzNB44tc77rB
MdfwSwnhojFdHcaC7AQu6PhY8LzKcCjO1n6Z/9VLMXvqg59Z6WUmlGd51tyI4HbZqTk13I4BYQLF
cdjrbBePha6rDKIGQ3zO9KrPyfguNc4T+jKLmXiFB+ctnn9IaVfpdQnmhGxmrkAvoXAynjIz7pOl
bcSJA784u2BEKZ8OGKpa7V7Y/Na7UnWyCKTGHqsInqN4i4glskT05/svKrsTjU2QzBuRtweNVYyp
qV/7X5u0wv8X5/0ckXgN8IJr+P9+vZM6IolWq5SoLO6H2SEu9aTTRrncq3g7MkIHBSeK1kQIxQRg
HD72HpFQFh/L80BxUqpoNvPt0Al5vE8I0ZMFzBUt3seTjBhVQVMHRerDXmLpX2OmWjAewu+/8R1+
iuN5Bsw5uf07GOW94YxFsG31VOU1+6QB0eHda28kpwq1EbN6TLy0mDYYEViSCzLpemEb9WE9Ldi4
eqX4+Vd+2VcXnti3nG/d8ZfaTc7B7O5y8Q0NdB+whR+y7U0sNO85hTRTWEeOWSOp5cTxp1EhacAj
H147X7C1ns0V2rsCB5KTKMM2k780xGDyxTitpAO4fertT/Xppm7kNcBA5SyeYTXNtLiDflL9eHeC
Ts/t/O+hbVPUHkqZJhK0k4TeT8xtPQeE5PJb5eznKNdzbUM5LdJavsa5FHyN7lhZjk0vwoPVN/08
7U681cd4sGPCHnMmLTMFCe8tvPFp3Guijrf/z7GLPa8qa81HOqhbtlnIQoOdvgZMnVya/d3KGJBu
zb6SiCtbO/zY0RtUtRFsLXVenRUo4rNCStqLDAx6W5MIVa8rIzHiyOT8jDlHtsLxtx4XViklwgLW
wZ4o3Ii2v5V5I75zujtKYTpeHqbEyRAKsb+0CeDcbW+ZjfsiuLoOk/lyDAz2pq2ky+egEPS1Cs+W
PkTJos48ocHFY790kDJLfFsIoGL89Z6pKmEHJaLTUauTy1XwXBhK2FrsdAZqZcJnmXEuAgoMiA3L
VUn/SSN7QBHGGGxzxMh3AuiV3wPxt4CpuNhS+Bkrs+dAaq6tegJPZKGvBQiIl0xB25lAgG4DDCYj
eDvzsUzrqk/74kHjci7Bpb1uBQAdK6+iAfMk1sNhGapOX5p9bTCLggeJk7nisZJ/GQG6Xrkf/3tR
0LHJwcLEtlfPNXWTwOyvlLCMrBPJvo51RV4/zhgFJTzFTP24k0VhP6xMPxFAQiY+fHVKwA7FIzMm
6YCq0n9cJrcO7TnFC2lj1MfGegtZtj6O4ewYqtu576ufy70cjVE59pOQYjn2PK4DtrJ05GdGY16M
6GHAWm81nVl/7agIw2z+06YmKkVumTjO4dK6ejwLufo0Hhvx2694+n7iCmarX7q68FNEws0KLj6a
d9SaopPB5L49//pkTEIXdOn/DDiYMYmOLtcZA3BWPp1wOSX7K5/bYhX8DkndPm3clRR5ddDM5ONS
y+J7gvtkWXd1f0Xy9rZCVgXX0/qDw6Rr//8ydsO4FE6esG4QG1lvxhbOkCAxk2mfEwPhOCoO8CKx
X66D1gxfOFJ7ioJ8ZrTGUMQbwOyf9+7zZAdUvSCWA37QaExeSUSxn9ld35CZd0V0rQ6tlcbfdlxi
BILV+1Tuhv5T14MZh+k5hVirBA26HRXAI6WcUjbgNuc85silS8i461B0iOvAUDMCsiODA9DUTT6x
jVBoTp9NQdUq4FeewIYLdwMBG2YdC6nOKMzfQzY3JGGJ1Y8lkDqz9TchqAre4P5hj3vlBlSVrKzu
4b8dP9kjShd3rUGT9Sen4Zvwx8wMQqDzBLEXkSL4mgQq3R/NKoRsfCay5TQnOX8DVQu6p7gsbsvH
IJR2zGPaHZ3rXXnziuomBc8xyrGoInSWoGKLSdhpmk1+Kz4X98W27YVJ1wwYsoXH6upalgQcqKA6
NS8nnzjsU1E45vj+XrdGXM+CduTpF6QX5KbDg7LvAFWNA9aJ9IEMzIhos6pChaIgM7NeFITxKZpq
USCWo9MgEgpLfWcGCZlGbxPfNFNO/8MKXD2mvPpZfJXZkgT0YHoBY0+x/6HOpytDykKBRFiVj0n1
R5STew3xCxQZsGs3bdF1JRMcFu9cCHUuWi+4xr6VG4+KcvzRs6gN0ve2p0yybsPdh/2a/JszQmSO
QintdfaBGnTVw0FP47gY2vmJPDO8beV2EzLAmKZ/qiF7sY9aM5N+CilNuSP7FedUZyQmWK73IWec
GiLFeGX1PeH5+9HAjqXeQ/dQVUIgQBBwUv1yGgb01yjr/UekXUSPOYNE6oLaK5q+tfVWHkgPX3+O
hSaBX8qp8zBs31A07hzN09VflAzUsGf9VDcNyIQsTod5HyGZonIMmG3ptVvmZ8dbtLj8wdSyqo2X
vOMgBvNFSF9Gl2AZXVDuYpg0nhi4ODMa4Jw5Ue8QyNGW3fs5TPUJSGaPA0U9Zeek+PVpLuiAqOgw
rDJBBCwxBtpX/KQkWIoOF7sHR2GBJobnEG6lz7pMKEZegNdO6pBSZpxaPpqMC0hJev36IZO/gi7J
6v0oP4eCkxiSSkchqTsL3i5INCvaf8YPzMVYJ9dFv0+LyGglFN3iOkDR5bY5ZNnaxfRcMSX8r5rv
FPp/8IeVr+DruV8fTcaJW9Y+/WvtKPglrx8hC67Nc8pHTKQkKRD+aFCmDiC6/rwHZWk8BA6pJTm7
3r2ZpMb3n1BW2EYVv0Vi6rAinNrPrdH5rWLThCBfuc+f2KG18pXk4JU6MkdGnFLS+iUKRfypQ1I+
9tOEtyMPOKycnovMIErKzzc0io9a5Q4RAS+Q+i9N6tqoA1tc8ieYIPRBHjCRxd6EJWVhWM26HgFx
tKCj4UTP2BAUm1WFUqVDE6gl6qXxn6fQZx1SukGEbm80iodhUke3H+6u46/MG9+qc2mocTDd6d+F
3j61U4Ax2LzMtt8F9ytFiPiLGkc4Ng9fcDX9SvMYE/oCGLkCTIPIs9dBVhP5vMZlad2RudjEltJo
QLfOYxRIJYVe6hDk+AtDdSIeUQpVdMG4JX3x2CoKzgsQxni2Z9UtZpR80kh8SXP6klWU18sFuWKS
eOV1ZXrbdvmAHYD5w1q8WUFzWtytKBvUcNI60BX4gTsVopeq7fjyy4CBHlmGz68BFUQWufIK02TX
RaVU/Qh2bDExGCHo0uV2XlUd/tEJ5BNA4GTi2bAexBcYrq2UgUOcuLuLaICGoOOYUYRC5xJjjXXE
bFLnk8+IQZ/JEUtwosnUKgJyLSsOCx/b1rtaztMqH6MEOa1f8zeeJQxA8H0Reaj+PKRuggGMZUtg
mcGsE5RpZDvQfOYH2j0O3xLry9dMSVeJLJqTXSulnPxCCjiUHlCQtHR3l3TKGoSrplDJmxfVaQtO
K0dHfRwVBp46wiqI5BNG7PBEH0PEqCUhd0wpE9uBMbYbpZcVgl1KIFyzSRiE9XUP0FrxlFP+CY/d
iF3ABx1fUST1LDISeEMYumUhcHqeFn4Fp1XHYGFu6x+KE9s4CkAewNNUidFFovE7vH2AjxJRlE5b
NUdb6hgN9OoQAW9r+j3EJermV67iocPHzMJfpP+Gl4DgjqiyZNi9C5NX7sjJqMb02VayUn4UaDB1
6kZZvbGeJ1KcBD1P/5mhoirJtfJJQ1RoU8o+vAmfNX3BUpMcenBGV3oNNaCvUGUC5UriGhDX4pZ/
w3Wc2RFVTSuO6L/swsMIZoM8Q68vJobmljutbCwfutnf1Cn5CcdCG+Ntj3+4Pj93K9HsRcAVDccF
WUxyP5mmcsDBxtjFx1JyahqlB5UYuaHKjpLS4ZgqgeMs0KX0PB7PZxuF0Hbqsiz2ZBocQoxGwIqA
SPDfHdl0a8OQklHcpa+qoPQwDtC18WlnfHG7HdU6tFgEdV8glyqsTF9MsDLNuCK021kojW43NQAe
YTvG1ArdM64u0KjWbXwly5AqT0qw20PozM9vQmf8SzXtfL/YSiLG4LLNLiseteZBC50MUBDW3Q7Y
d53La2nO8mLfRSTyDZ9eIfQyZtcr0ihuqE6T1W6cZM7E+HE/QR6cmrrrdvs05Q4bPuix/rKmDXEE
872dqyRoz3bFUlWtTUHhKnGKxNEx2zov1s1S5RR6qO9Z2CwXvQYZgdbxn5AVe3OnCaecut1CaxMV
VMPchxf5sl/CpDpJ2jHnuiULet1JSu8drqNezE8voPI1ENM26ZY9GwrQQOWsqUsCLdlOD/tg35fA
LNcYwtsFv6Uznr0JKX/LO4G2bXPaWRv5RWtV2nBJ1GV4NXhKNhYENoKSQWtesP7Dhr0NZDV3UIDV
8otLpAjtjBj9fi2E02dCJdfXSh+iXOOHjfiXA6UZskVEt9d2v2QhB72kgwkaMrSTlQm/uwoYF9CG
OEuRsHEIbgTxTvDEVHGw3w6Q5aP8SE9kRPuswKJ/wAMJIWAOiGTT2nvQTwvuVxghBXdrtJvX/8Tx
ZEfKms5affH7O1A+FkipK600aaYWueAEKTObIwNER9WPcTeIobYVwpsHKF7i+6Ou7VopR4yn32Ep
W+8/niSGcVUhNqOS7s778jCKYTA7jEJGD/XVQ1JL5e+z9cxyLh+LHK6Y2jzS1dQJJAPEfhYgHlqm
JY7e/Wwx88Oa0DrwMPNb/eIPsqVnwwGShEnvr27gGw1zFzZU03Rbbb2Ma1FGJKPvQ1b5lO4SSMMn
QLzmVSvpHusu9LluW2Tj7vCpYe+hmv6gHEvhPigVHgrJjThAImyOF8rLAYIpeGbWcYLsGSMINjLe
Cr3JMhd1Z25um++ZNCSWIqoG8ci6ynVCcvc3XXtzCVntfda6o13UA+HtGzqC9J1/E7jeVmsTfbMi
NpjLkf+hNi/8kTezjK96cBfneYmqpXrX1j7kYtu/FOOLLeV2TZtOkKKq48GcbbTq3Enn5Lt/U1MJ
x0UsMEIG+hVMa/SaAFLyJGGtldSPF7E6OPCXJv468KN2Bw6KcM22gkmyCieIJBMGWW5F+oG2ZMue
jcv6CVfR8d7ELWo+ikc4yXleXKs79e1zdDSBrgHN8L2Tbm+MhL1qVpvDics0RBnimCsNoTBrT792
GcG0VTnDXgylc9SW93jfhh/9orYYK6MzDFKp8XnFpQwTFBaqD9nW96KMegr5Sr9SF1yUCwhKQiim
8eP2w25trK9DG4L0uJ2wmbwTKcSkXfzS6SV60SoCcdYSqPIFjw+eyYM0l6NGe2NrTgIMLyE1Ywpe
lKBhdNVCXa2V7UObxlJxU4fI68bvDh5TroksY43tM1B5MMiB/CMOnTJtfgBYjYvDr3wy3hO7+JiV
BypUEMglah+n1xvxBedSQmIydk0sEUXbNJe6upLSAd3T3PNZQWB0kJ52jXP9lrMaPioqT6UIp/xF
XdaGmydkyTCZjKolO0ROtbC9UynAt4vA1Ud4yWtEGtd531tQfMgaRI/laHFue6exH4BJfm3c30Xy
7ZIaTNRl2GFe9VLKe+vMMMMUNyt5XGt7EY5qdx8v0kKsYo2bV1hckrl91zHFcnHCo40HH0Fjh4mV
fswdmsqqZM4aX57lcW6arYBRfNQM2OsazoaxP0U2AVPun/CVHVfdf/ieeLCeDgtYCtcg75CkxNKH
TesQfCn+g/jCKJeXVtSw6iqtwMPxlMFcA8BWChOhg2Ha5akH9oCWgKepKOJB62Yb2jhEB9GxQ4wk
a578dXQJyt6lQZMuyRMXk/rIUmScHRenWP33kaD9MMVjNykBkNnrQZ3Us+PABdiqVPpcJvSZsMox
XTQCbaTt0oMwz8Smp0buTSLmbClEx2sQkFUUbHjBjhvMya8dP+kFdDCjCAgX537GJ/9Tdok0XurK
AJkZhYIYX/SWQTX1ugSY0fMN+bwEZMe44uQ4ohhLHthGd87dWmnIunKTy8I7oKbr34jg1BWwwfed
J+zND6h0qgmPa/xKE0OHJrNMo10eMHch0ymy1OdgTCWy55JdRG4sVc+liMKNNrNQxXniXfULehXV
Qmxk7rc9WNmpjGRNtCFN5OzWLvMn88yixiNFukq6Ofm2wrYVfMyBtawrJng2SBJggHpNTIOhnq8k
StKSoY69iU3EBNxnYKhNwysbPx/Zv6UbMtVJDd2IZ+Ii5KVONvPiIzp9zEX9dTTFG/rsbR8HVyIv
mn+XzPMgvb7cbt3qNmIlzjAy6jlDOlG+4Xgk+4PEANZ8r7wZLudhShACcq6jgyt9te0NsLFmTabB
1SVSTDtwysMtyo1gPuYb2EGp+IHxIfkCdWayVTNJvRCR6V5KoHEBdKCQwwfiv6px6MtlG4TgUUvE
VaOH+IrgHcFGCSvCOyiEMFuGRJsHyNV/VQgm0Kyoo+B5B0+Ok/BvBlzJvhYJYttcGnaf+e1iHy8R
I2WoEMBoZFdh3qXaAPEAimEiYoNNR+0aScKLBZGsOJhyASvyyVTQJJo1vlhOZTjjwnrmQ0iXU7jD
4jr+bKNE/BZ5O504lLFq1JHR6pHYdqGYLKPpfpgs+WKcg2rrygQGu7+/K6wBApGZS8o1lz3cHV/o
cHQ33RNMfHyAC9PoJ+2jW5ZBjhIMOk3mqqtIDD//CgujYO2irM/3jeMZl/6K1BLOv6RYXTROiYze
uqvG6Waqity2MQjMW6z4KpFUjuKCyw10xf2U4MOU269Rng3RARlk6ru5UxeELiV9li6o2YB7Tl0g
m4N2wnQvM8UxYkboLJSSiVXjGeoYQj4btMU9TWUsYvk80b30HSvTMNO5E3aqqDQvxAXRMR5PdhP6
MZBhcu+ODGIX9cVsm5/Dpi9xbd8twY2UmYhdc/AsZccpJmVfKt77reSWLk5NWoFbl4HEg6pxps/K
gZBXjZfrpymwNA2kTRnSYwX+6bKxILD28Dp4Y2KUJ+WhcUCcy/R/FIPpHd5KcYe9A+N93+02eF44
5yndtnhjVRDYlF65TSrq4jsxNPva2L5cVLLyt2XYgH27dKfnT5sLOp/dbmkP8kFqhoVWrwubTHfl
ZFD4Aoyl0AvdHlF6TWuEXp2Eme9POEYh7yTOYDNOCd5Iiv1gYW9hXWfCUkJIvf+vWOEZ6k4622ax
dv34UKkkrPKcfmBz1kyI+aNoJQcfH7wS7sfYPS+pbdazFURZN8uNf6qEuiZFrG38WoY0vgam+7ZI
wC5HknnXCKEtiX5JaZm2yhZo5r9BBbI1ivAQ3p/WW/qqIBiw8hL3DUvsXmQMi8refWZaocUFJ1+0
B2BekODEmKuN9wCPfcOhHWdpKAiVegC/3zz98jjx3PCRA/PBZIcHyO1EJyDwrSyeIbVyHG48D2B/
boT3yQp8QazzPyE7Td1L5B0DsXP5n8eSJL4gxIcre0mi0eHV+5lcmfFefHrhLqNl3dqPPc8AXSgc
r32gXUWnUZSDW30Ylo6daIdHwEIpDYi0lvgK8udsZwyJ+wXIm6YjU+2blJUaSwz9XmOx3Xjc7oYa
CjNR2tBkl+SyB+RqxdkIBNyVhIhqG8YG5Rp0ADl0lT0r/c5Eh+7BHuP/xa3qvdCqd62IQOWqmBvK
pDzmdkfglTKb60wkvbxYNvQ0jw7EMuYm1GZ55r/aGoXCA1iR32HhUmzLubyvOtACikE7Ij3ZZU4y
v0F4kHhMxCQmQCn/84mXTb4jUGpTO01wfuGnpGiDdWJjuJEr+Qs1gp4nieAiQGlTM1zcjrTn8XoD
LAkZD36sl5hREjgApd5PPTT/i7BRYQQ7n+E3EL9oEs8XTWdmk0OsClJN4nKxX2Fr7hYntJRErTx3
HLyNOnY0XYpKTBVYItl4vMcdFhsRb10/AzVcqFIflOOAxI/dvm+L+rbaAKsH9CJ7TcweV4KhLRlN
NJwSyzPQx2OTVno3XIJszB0Qfz1UdowpKFaxq18rW8jpqRZiA36KSX2A95L9eu7ElsYoUDSKGAY8
nPRRLbmsScTXLLmDPOgOyETIL6Wn/kgcEu8KA9lMT3on+aEnH0uFJqhL/RUFFp3K2c+GA7pfhyWW
KdesGV0svAJ+yYGL0FAJX9zC7cpbppGBjyZap9nvjpfMsvx1gNbLC9Akn5C8jKVXkE9ESRqrESBl
M5Gxg1EiNrTUEQ+kK0lqGS8VdyqTNrc4lP28/AP4R1CA0nMUQIxpMfw6SVAr/Az10cMD26J1Vk/k
ruG8b9eyCzMOoU9bfBR1xn0AiTVs9LiYeCwxVTUtgZnaEIs3dyWW64MEZ9BtQhZkmTCFyeZ5Bc8M
4v4VeL77WZ2FUmfy9IlZdLyDp3p0sS1+yXa/U3e37psiLg3QxNUstgvRpOBv5FKVCg7363uxFMYM
A9ZnTGPb9kuagohlN3x9z7dat3My9BoVUFgbotKv7zRERLd1FpI8/ImhvSgea3+LXPtcmi5I5YKP
vQ+k5MQS7ntLqNY9M4wIOLVW0HIg6moZjqLXNwskOybLl2fBS6HQ86SL+nzk/gaXPc5TyRR+r5oU
KQg8J5x1mxzc+BRwJCK70+4aDgdJLVio/I7uLL3M+8QZ/u+m6cLOiIX7NZ7k8kVV8QLs+8Wp1Yxp
3DPnPy2cRM5Ed191kAF7hNAttne7t05dK/THoZBwOIf7Vt4p6Xl6F/IKbMu6eaqFd1VCjW0QyVXB
SfRRgRhcz/PaJyJe/l7PtT7zpCO3U6avt9DvrjajBHE3/2MzzcaaJVGwAzWm6l71V2dqFFMu43hu
BwMhmY1/V25Esf6xYyPELv44lJ/VNijdXk2nSLmHWgLv7kMAA5fza1Ts1UGlMLita8ElBtMeU4gI
0AnI7KdwrGRe7O3AQGMaoyzKkkWVDCtuTWivMLQOq49EuUtoUU4HqpjUjbF//VJJ6dK3DvuKZ9JS
VU23YsIADRwK8Y0fPlR48ZZbS6XSn+m4yu03PZMhhrLY89vfvmJohaVtfObb5BACE3zAjON+8pPB
1IGHIeLnVP20IrClnFFZvxKzfx/LxqZ5ttdi4BuvsMg1DLe0t7YuMvTQDNPAig3Ycz0bk6IDd9EK
52z/J6PNoDsWDqQRiqUVLN7zHMvglbnaBBFgOiJEL3P5gkYiObCCb3U8tRQ5JfARRG8jAwu3e/RR
56/WQ0PpQugra14LSUZWO6wbxiRqA4+K4i1nJhYk50RJ085/FXjAKjmG2a82irpGG/hm9VVFxgg8
WY50jkdfLFkirWhp0dW9wr+UFbmm7lLQ9R93zaM6EOYPG3P6FErhdSsMX+vZvXNSyDIkMSz60Rme
dBSUrUtgYTU1YzLHf6XIEvkgspabVkyty0AR3KwWuYEQlMhDetMpe2AJRsAS0uislFESgRKgIGJq
1xLmay1mDxi4X6jt5QQsvI6UbN6widpDsqIRSe+ivhCQ/EmqY9IZCH6d+N5+Br0VSWpfioqUDjxf
qV2a7A/Pci2db8sMOtWBKoYIUYkA/uZ4dR3Pwgj/OOaoOyVNHUeVh6foNq7VadhqVl9IT+kjzS+a
P1LLEv4OO0jrJDhovpa5SpHVHuCDCgtIPxh6oL1DWB+/ArAgkPurS4mkGGFZArt9z5c7iZmAiN2v
O2VFW5ab1MeVeQ7V+5qn7ut3/CUKRZV6zJajix6bKpSpT7ddVUgFMyOiNE0Qbkg4Hv296RDLr7jp
Cpom36DKOQpNFCkzN7pc8/+861pueFwhynIn4i7zIpdFHgxMyzEXYag0OlZRj4LboJFGNngDGV7T
q/vTYqa3J6+4wxOImtZ5c7k/FP7oUz3pR4hccTjxfwoaTeQbBy2MxUOewW4jp/bK2Bb0m4jvraNT
9l5jjUgz+43EL7UOrPTzJHI2lkXyCtJjoeKwSZcZjLwpn0WjRqaN+nKh2s1sHlQXn0e2YozodqJe
41Z7SJx88RQSc3b2QYRWdPpW82vOhBYvdOewEolM+4wnqi0pKp/sjsyDolTHhi2wrnJLZCDK1ac+
M4pFNTfhh2bpSFUxrM7Mhg4Mg6Yqkuv6TXw1PYH2/qTq+WfQwhu3xxNWGHdGDQErt8NJuUHUzv1J
r7CaH52XhxQWH6Wq6VTDEbV8BJrBAwJ/IStF8d7HHIOd6qbfY6laR8G7dlsYrt2q+P0n+4CS2crG
IPDDdlU/Or3JitzSoA2xwTy0mwPETiz2zV7xeMQpJpoyfT3byMJdz7uCpq+3ZAAOuraBNdciy1R4
UwuW1xsubz8ySMnHxRhT7XakQazApJu5oC7gpc8uj2wBUw3Mo71e2JVaSVnUV4AKB/CwfKKElqQK
DP3XfXRRs0yimcwF30avVfIESbqysilXV/8HOMzXDf77fpF8e2Lyf39VzQIVrWB2Wha3RBLmoNg6
4SQw5Tx91QyEUWZ5m31mqJivINWZozjDbMOdc2pwajfYW5PRV6LVBtgylJmsV6QEMWZzBcvcNjTQ
H10gq98Xblp9CRvURbL50kn17HvEpu0I3KJy+4AMtTIFNzSWAoSlkvAyonH8zu1mbhT6G+kNC7WD
8kLoxxWB4hH7GUXGA9wykQpAA3i3++pcE453Ax1LT+l/mcyibb8HLM0YUkWHZnWardcVdzz3jYSE
gxwWtzS+7nAE17WIdEWeGxDflNLKOFA/Xnjd3tWVabU7Lr+JBgtV9YITpeOVS/F1DnsQkndT4Vd3
rX43SwiFirnyQ0uTiijonDgzAlQ6ePTj8ehPVF84L8R6q5lQ/zPd/zOPNaFXH1UJeQb6ecQw2s9B
u6+VmgnXITytj+tnNE2JFDOlwMSyJ1x8w5FCZsvvPQhmHSBZjef0dktePnSMyERRCCvHs6ugJ8Wu
hLyQL/Gg345EegBZQ9g+hNhV+coLMqxd0/iJhPo4t5xvNCeKwrONEl/U/NF3WABwlreocHEj0URy
sX2MA3nwfxygOTT2l5bpcXwdgL7V6sPOgOi2EO08fKInrFOAx/cL7jchcMmRcHvh9ym75k6Dl6xE
RFwMS7Qxv9yNm3oOqg/eRqNkjHeulrmaMGSRvk59MHUW5UuGZNL7OvnaSLLm1QikSzG/avNtzUzN
F/AHjfPHhQYMJXAe3rPo5eyFcinPSfIJCX3NWRQugFso9Sd64vkiCxeB62FZY5E+dW0cg5cucmB/
LRS82f3OCqDc2BPlgWSzKT/mqYBhETRpB/12YKhJsO5ZTFNiClG25QUBVq0dCaP4v5QpICsXEsNF
ZoGAe43ac2g6pHY0Ce/Qa5mdJMGLxuuw1n/K71gthCURgcq1U4GqyIJ3DCx9JL2h9UWdGoUNZf4K
LWioK8QJIvYdl7+yG9cvtSmcb2WEP7ALlBv5nG9WSn25OJt2AaRW+1w9ZR6VcTyG2lioRTKoIRWr
nXUq+7ZLehCsySSJxKnC0pJqTs8O3rOQ2YPALBhbdAvieNSPh6C/YnotwObXfasfRcQtV4PE3sFM
x4djBTV8GuNYiJ/sCmJ83uIWB/Qt7BCi4qGwAxpZexeSBZApxEO8DlcXW250ydIkaF34lA22md6T
C8or7v2zXp4SD2SX7iT+liixtMSD4zcnH05x4EBCbE32ZXZWv4M7/Y0P3f4Qwzse2TTCjt6J+DDN
bvYlp8XmWCLBExheAsTr6aEhEwUrhgdL97u2th0dLnIKRCXPjVQ559WGD1eQxK0bWDHkGwWvJ7kJ
HW075dy8owRApjFrjjqYeW/5Myl543ViQXADbxay4IFqazUW9WAIvGmS/hg1jbzjRkw73CgzoDN3
SgOy2AtaDQFadtUI1+ttE4mjW3igZfE1HZYRhd/ZQPB8iGLC3p2poVnWWaCL181u2wFCPFDIt2Tn
rqltXlKRYZsmTtDJWqn4hXfRrFLCbs3G2p8S9NtwV+TCLsP32y4WMNfXE4k34PnXTGdti41fQsS9
cn1KNrsbdTDFXNrGfJZoYJ3gKzCxH3bJB+bqIX0ZDkd/04qhSo0/AInEabF8LF3z5CV3cCHfSzbx
9rUnvFyvv1WDFrEZmappS5/5+mrCFSqB7GZFzoNNimCD4tziTEAkzH0fE+2tXPisSTrrmpEYc8S9
Ik/MjbpEvKdmhXf16v7LC142SGK3akVxcdppHmdHREa+fhgoQnYKgleMO9GQ1xgOd3yrwuzLVbOy
wzTybVtPjre3c24WNkgU1MCg9P1AxBQVgKq9Kqcs2r5Y/cEKsW8FGvRfpqecfiZiJykLs/WJAVkx
M/LnJyeGNDScjL54GWNLAPGExZFhg05hJNNaB0mlxVW6bq/iRNQgi1KWC1CMaiil1lat/b+3MGwK
p78UHasdxWUX/v170sTQlClBTuMJfv1I5XvjXxRr8FEQQ6CXQ8dZEXyiErVDPapEUlGMUkNHiRB8
iijxP44PqTuR/fbknQUfoh/By7tU6iB0UnEeqNFAqskWCKui1rw42Zg7AWjsDb6JoiAfBNWQnl9x
cK2XrazBwkT+r93eXnXanIZb4BOVXXNauHkRReQJRoSKOZneqUWqWyVkF85kOPLfeymEvWo5H+5U
t1VKikixPh5Al1TymFtJl6PcfOKiRpP35evw5SvBqJkIp8VJTjDDFrUPg5IPSw3lpppYmO1MBmz4
bxoXZGw8LbcXVSYu4Wg7luhKONCenKI7nspTUJo2+lEv16XuQZTTABk8HaWJm7gtPxAvs+l+5D2P
9MyEZW6WmiyPkshQv1xioDTzTZRgJa85/pCcJfKG6WKUagdTQWkDln9dYzC0bPYCdoYQ1S0SAsaE
Z80v1Dlv22EIP5Qgyt54lv0QxL7L/7RPIv6NaU5zqEUz+Hyx4JO/9U3Vx65uD+vTDxGpgGBFL3XK
Hkh4KUtYtUkzEb2QmflQnF77BEi2/ToNcG0xouLmTfuuobuETvdL4hlrBv/op18K6pSYjlO+TDLR
LryKxOGci8CeqXyg0xcFXae4lq/GnITQWkx5EDGlbHOEnMmQdQ2zcBonMKetzBmYYiw7p4LQhZUO
+kmTfZKkks2wJPcFvFH8jsQ1ChwS0cyvQqrwnbxB/OPblFnfjyTzGoyWOCZFtiZj5/qYUDAT9usJ
WO6cE0PERsAys1ruPAaJrMh+vb+oF7PtGPMQY8ifQjaQyoky6C6MqW40PLfmhIgD20tCdS12Vvbd
YalUieBE2QLoj9QGNM+HAXrQ9+U879+d+DzbydsBZSMFlJZT3zN/GOHJeZYuGA75eJJweZMLuIdX
lkug7UP3oWAB8NY4F22by6rYh+lNUxC2xCSMW1JGZ0M++JFsbn/LjmfO21CaYV8F0lbq3bjuawfJ
djlgLxHLb0sTPNJ6rHGVzPedjqwWKMILtZCbJ/y8wJpJtVa3439fGRy6KSoEuBWI4VDxKPJA4AWp
vfbf0tHbzJouOQKycaT+wGha3JrgMoDHbgdK1YS8pCryDOX/fPQWrOmH1lH7DsUP81WYKQDCy6ld
EwvE1X25JghHFlAhmALaTYJbki+8/BS5sW2iiaNeORD7MPoKOgLxjngxuzBYZnzG7/dlNXZ51zxm
9tgZ6OYWZhKa1rDBEAd30jHY8E6SucqV+9NGvnE+14IgC0Yl84RMcA+NPkejLgC1ti8BWuWJmk/n
TDrVf852plsRrbWjruwvl5ajNSS61IzH08YK/GP7fWrBmnroSuwelUzo8SSZtjRPBkxho1QHKHwS
P8aiBWRnKf6kOots+2n0aCWDgNKWABuspA45Dy711SCuiZJjvv0JxvLRXhuXt6jx2azyLCSv8Xnk
PpS+0ZWdI1cTkREJijrJ6I8lcLzu/yultLFihCddNooQHurZe7qU7N8O8DkhTqVbKgmxnaHrmA/W
9S0fzUfarUqR/b6V+YDNevQWOr/I70dR/FEgMz+QwkFaat6r2ZeHu9yhPLiKqUJlvQYD/Plm6L43
JJzfqVvmYMxri6vRMUIrBG/6ZJd6MpGQKTs2H3tg3+3Nq+LVUQHEsJVGJBj1OPDyiLEHuxR8eqQ5
oPPnyTRAO97SR81Des9iq9uMcTQrz0gWqynfiendVJrJpTxVkRd3XnO2ZTnYvmppFaPFQxEVBmhw
JAHu7CBb0eDJg5W0kwvTmAx69zC2fejCYbFoBTXGkl9DLO+o6eCx4kPQbD5xssIIVNkp45U3MXLq
TUTWeAIwSS+j1jw94d2hVK1Swp2845/bN4+f4s8uRosoBqY19RPp80YzD1ClSgFgm5Ol/hLoV2j8
El6Qze3zzYLu+8YW5aWYX4yKRhX7dysd7v4cz5VvN3+I0eXaWsNycYPpfAUQY12j4IExU3dUmEXA
Uhfe1pAXQtUEcvHo34SyKkDY3BqeRGKSiXLfOpWbBdkDaBxGK1cOggymK95tNMPdoDE3QNbpt/cM
9JE7WfIFvHcGY+RN7Ms0j/MsqnTeyvo76diB0KPSQhZt6u47uvXSO8MeXjAclySgZVzkH3bphJ+N
ohpPuMiSjch5y7UQXx5O6nPUauASiU062e0ihuHU5MC5aPe6QGCmx68CKeDgz9p7BZGmWI9ZtJC7
r7HnyAaHqDBflPMVcbPqhun68xW/g37z4q1sVDQ+y1ymNWqlGtbTnN95HPub6OPI9hZmc+KS9K9K
NyKJ2pQ4B3QI3fxBSZwvfFJDhpZMIQnJSOSBHTrUCjnaEnWayb+iEHvfzUYs2uzXkv7eBabbR79A
QDrLUJKZo7LH+4IBs/fLq36csxfQ9pcvhJlF4xF5lj5o9Qw1N0CY0SbBzzcY7m2GZLelb/Gz4sFF
LUdFLlGnn5J8rFrUmVnOL0YdZZA9IqTnT8KqLwSst7n6yu9djxgkm6x/mUxT8+0iokKZftNTjxo8
gZEkRD6rrqDSlWlegWCCczjxc/LNzWTGpqD1mj/oCiyAKmPVP9QhMgmAfk4K4VcZ02BEjblduRVo
rIw+q4pY/TnFixBLOrfjrDzxptEHz/vKEdS24iUJejQxXhdQKBZhB0kGhy6wfEbsE5rWDCP0QBoi
iJoAapA2TdIo29PBICqCvrJ3XGslWQc0aQVzggkYYMGCvwLZ3wdWOy+1kHhkyggwxowPSHqOvwhl
yGIGzki3lwVWY9vzep6gLyyhQTfR8oEPbX0/rqdO8pawTYn9wgCMCOZnGyng2VEh5U9pvIXedBvZ
8nD+V7686GOadAvJfq6zKhCWUFEXQiP2Q3hQUJf2p/26DP63koaNsK9ez5a55ZF3b41cnH7X35tx
x+QESmvWCJtKvkrbpbiC9bikM0KGMftsDdp5CpsC4P1o68PPZW+yuxaLvSUYxGn+5Wp9GBzMfK9W
68SFnk/sWCZqNlEbbnia3IfSh2/G4BrPWbp1SUaCoLsW362W1heTJGueB2KWtNtFhSGm2Pt+rkpF
cWJAM88pYXN71eZLsk3bl+Af6Fj1g7ELeBukjBPgubIggbuWjoNI62i6Jh4DkteIvNh8xfrzDjq9
rHDklLiJjm78efv17354+M+wVA3X67avqO1wFEnGmyctfRNFFeMB66TFr8ZNG7dmDcssP/qdF6n0
GWvOiM+LUFo03dQmrOdM2uPHobYoSXr3d5DWEjB5Y+3S8fn95K59ChQwPYWVvP4SEnYkyqKYzM68
XcjUfvByCD6rbt2uTJt85a1h+WrMSp4K26IK+jUMcvtgcacOSf8Os/7SOOr7mPZryh55h9pl485e
Ub99m+4KuS77YDvzmu5nj0IB0et/1/8IgabI076UsNYAhafHw7CbtJf6tej0QT7enZJo9tbyUuuI
NOpm+u1i9y9M3OJe+psovTtd7UjDrbouwDb0n48DTzd1YgizdMcFUjd7HZkri6d/dJs0j0pXpD7D
89Q6JkK6+QcVJjjrSB3eI0UqsbRIWgBrPBprqdIdmT1U1PN4ikfzp6f8ZWoCKg1woQazz1nkkEqv
+PbOuuMX8ohNLMSP/wKK9kEJF9RyODo7Lz2Em+N+mZQjnPx0eh2yiXvXNJj7nmDVP492E2EhFm+U
i1yy0Ao8ozW/3nWfL+T3eeYZR0dqoYIQFl4EBrdFC4BMd2/x3njqriq11kZR0QCBSo68QV5LcDzb
XI32ogn8qNKG0aru/Y3K3lAOITJbgQ3SgkXcV9X85oO5q9PaHofZelcYM3oI3fwqneWFJYNhygmA
4ZnQx28tuOw3C8vrXVc396fEo3H8Mn88LAzVlqkz4AeL7wPeJTfKAmxNts9D4Ogr3d7xkcaei7qu
cyKq1ptAhbRWF9FIzIHJS79BLT+D+HddYbgQgrW/aGca1oZvPYMrXGDGtG5C8rzzVRK3SSH51JY3
OnP/KJ++K4MIXlo9VUTEkVEsImM8MmWfedLCvEQcvVbghG2OpaDBcHEw8V3qt9gi1RXTwaSqhDdZ
/OTM4qxkQMqizen7Z0etooBWajxSnar2dLN7T6kcMNN72W9c66U+VWCLSduW2OltFGYPjjw4qd2L
VMnpW47jwfje2TOBvSa6r3mVOSFabFAVtvEluPymTOn+G7iucStZM8Rk5nvfM7hPucJCHiAC/uL5
9LL5Xrt0j2rOSQJS+JLdPANgloRJ/ZLqdSZTI5YDO81Y8W7n6707dTM/VcEGdCDZaZCX0WYKTO7n
AG55Y0+22kIMBLN5ZkbPab5yWKW40iHd25vqxUAnoiOLwgRV0hf26rHVLppZiyFxwzw5wxD9811p
kvlP7w2Gq04cTPvKEi6LFEafJugQFO/fFiH6YNIWOq3IfqFrdQXBKdxkF8dm/jIkyt4ddw7qzrTZ
RN+RWx+aSvvEFNq1E5SGfa1DID4Kov02mqoYhvZzi82kiTbw6VdY/GsQ07t5Vc45KiEItgLYhq1F
BCcbXNCA5VT3p4L6M940pb0/e+hSp29iQSbkMaudYpobqhhZjUSd0tqAMz3k5vxG+eU1xCdQ3IEJ
PtjvoAd1cQImxAxkcW4FBr/tuAmoZA+LoDbSttiLW5EI3xShJBc4b7L4aZnD2Tpvx42rRQU/dZwQ
Ppbwiw23tuq/SeEfibLGLBYkgGzSylIWM2HQZjcWI010KjeP7JNruCOyCd3kOJHc8bFkXcvRPR/o
2W9bXYtxpvAllUYP6KEGKKy60ORjRp7B8TcscXrJ+5xpy1ullZtSvKDluSxCF3xstheQqRzXoZXv
wQ54ynM0KB9irQv0vOFWrHm2PakJa89ILDBe35kb2moGhHY25rEHdnAmcohHmDOMLStlAXNad81a
nqzvuDHTR8mRgFXtrDVzrf/VbbAVRaqNFbjaM3UJFjRTBs6PyRKyCoHS8yHRBmhuUXjTkzEF2+iD
pap9j4metD8ZlzFNp3CxrzMm9bu6Iv87d6fQX6BgbfOzLy67EHp52XmUzopSaMJoXRoKW3HgcQQO
30JyRk3ofKNm1tF58IqM3TLF/9E4XJi5BpbEZkHGXuIora+Yox+99NDwGuMT2I08nJMs+Lkmmv3Q
eWajVmZFQJe4YEgALioGIfrwjDFW6BrO2GIXSMMOa4BtUmfaIk37Era6Fzmfl1Jj40359apmaLto
NmtlYYkRRHNEYVTkwBzG1emEvoid+JaGtw13x4eOwAsFw1PY/CQauLnzfdqYnrSlNT9xslztmV8f
q6M02+yJOqW/7x0xEjkEv1mu2TLcSZMzHKlSN8blmDOA+o3e9b36t1TcC25gSygF61rKl8m6p97d
O9u5mbJzjlRPQbtKZCvl5fUs+dSkLqsCdpxIRPdivWE+ygCdyXIA0FgZ2gbPdWVHeelwqxZGT1nB
IUK0UE922YpKBN4u5QhbFwGEgpi9X2IcBwbrNd8lQCBnKIppU73d4S864NGsWMxL+9FO5xmt6EXR
u7a7hLi1qMLbvkGO9iR8rurRyFNnXxmIEW7rTmQCsvwoeE4Sp53pLHOULL+3g/5CaWrD7/NCmlLZ
LbKSoThjaPfXMSLr6Tna+Q1rzpeR/blrYIcVQwXG
`protect end_protected
