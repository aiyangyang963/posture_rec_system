`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
EgsHeoOxdUxsX5gIKiaj0rabVidhYZrAC1ccO7uW1WWUY+5F26NMKfuRo2RbzpHAhKg6YWmehafX
vTPGaJRKHw==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Z34YzyhCkqWVBd+wfHLLkUW/H60lDZ7DBcaAzQK4qK/8LgoJdsH6DZ43BtKjfZhNz/T8CrFXpTq4
lXACmrJsvh8DNPmvB7LaQhnP9Q1UWB/2BUP3fAUHMA2d2pKOqEj3XF5pbikvIPiyQENN7Kn513bC
CvwAQIx2bzxkiYX1MZc=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
SSMUY5NrZw2M/7w7U4gsSjNRmWfRCxfALTKD8+8C1h91c8RWo9X4x7A5m9YG0Pa491k6Lxf7I0eD
goajxjfLKNI+buWpvfZlHEcU7678iPGqz4g94c5n80sa3TKcwpV6f+p7C93Rto4JgUHSigA3gLBN
DzpD+6xOS6P2mkrRsQs=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Tbb//X7l5IJljgHR/Q0swC7OpOr9LwQv6rxLgPXOMJNm5TebIkTTeQKZBlg96/x0gqqgFX19ZASr
qWxh3YL/aoYejZTUMHYF7ktggRgHydykFFfRo8xGrq33bJ1LOeuIQOZyZjZTB9zCoo8CMX8wCtcA
0ovBA4GCY5VFNLy/1whSrZs8R7CLSdrlxUJTTCXjF0f+Tf8OyjSS2VGyZfJbmSNnFJJuItoBbUO0
6qdcZfL3eQrA6y/AWPiFhGILWhBAvVGEahvuOHYDa8S1IUccHMOxQJtq0Y1UqRNB/qNmlHUKL/iH
IEr89vPUXnsfHTV4I+xFieSKz2LwzLXsAys4Yw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kfJNFYIhzZvlPwb4KI2aCH6Fx40tZkxF1Q5EfJSPdq2JohdV53Dn2x9HbgUIqvISu5UuFwT8R+oV
/B66+AOKivg+iSCvhh+HSv/oQNtgHeIG5xMgV8d3jXD9G4abV/g3jySuWrjXT9Z0IqvTQjqmKOR2
9nVDANRSJiSyM0Y275L4ylvrdjL8Yim0M/e9k+N+kNYfcQAzQYd/lfTmcdkn74/0qt030HQ2LxSy
A+NwqYXBuB4VkkCPvigd/s63XQNHxeHfRZs7q0iWos8Jgu9uI1zA6ZN4O4Cts2V9BF+SRqJdzrLy
1t5mzK/i0gmdsb8ds3y4b3AMet8PeT7w9sZc/A==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
MzDVqgEdc7DZdlm2cItrUQlry/9kVuVoApPpWX7zga11t+tLgAqain8Fhjl9Q1hFV6Rwv6WUUyOW
dL6uK1Pj4Tc0mqHyEMvAW2tHA/QcK0pphBofEd8Sd2oRBJ0l+XghTz/o5eIVzoxDF0h6fERIgAw6
PZK1iaI5d5osnKGqaJVhxQWf/M3XiOn9jCOGskyvtqNiiXNki/oAWPJNgm3Hb599C3ugMxNKGT5x
H76UXyZbcrmrFSkYz6XydewUEOb2eruDdZtf4QmJWyJ+WqAHgjSB7kcn3UfysW1iW59u7oxSpMgU
oLKWKFtXGSzN2+DVJ91qu7hIDmX5Q2X//JK4Cg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 296032)
`protect data_block
TFQ5w49J76k2LAtvA1zQhtkNO82XuTLgFS8rijDJto3TKxJWPfQ2k1Nnat9jk9idYEn3BCXTeWSW
iYsVvHwnj5tMfmP8Y5mub+t8YEwlmtbDlZVU6XIbD/dABoOkQ7/dRWsGY3BtHzylz/WwBsshGw/c
QNRdiqzPiCoHjSRXkLmpl4ZU5mQyuKdHm8u2JUtYwzuaJ/inKQkiU9bQAAIvHOsSMaR1mW4yF+v1
7hvSifS6PYCU5vot2RAyfc9XpbeR2sCezJBazlZzOkvdGIYaS9CTExVgTW8Btrh2X2rh+sbhfk7u
Qh6gB8n5nVB+TD/UBdVgJ8b/ADdqgJ53MhERpPZHuRaV3BdlofiJcvSG0Zh6S/lP1W/MyR3SA1bu
wts9TO7JCBq3UmruGBOCysVSdmr5XNyc3mKtVkT/QCxcFCPIujgMT9S4i2st5xUMJ21KyYWmpxob
Q9dYj1EfU+SGHJLhfmq64l08AgCB2O+TPeWwaX9Qk+8ZUS/EFzCL4FeS3vfffp5yuo+JjQF2WKz2
7VgueKCIkd9fH+gLBSvXgjkj5ZFR85rVEjAho0QRgsgKdYvYBn21iXnfnHbv0nNrXVf7ky9pEJKw
rIyBiow8QrPGOr2njQkSuvS+U4pnPJX4nQt//XaJ3Lz/42tZhtFC6QQQQIF41C+04GYlPcFZEoK1
B9WfILjUo3jENmeHh6A4YKrvLt1BjMLK8R9mBW3AMBqWJlYeK6BpI+PVJjZ9eAZxVnVWM5Z5Suy8
AGMqUvjqxN6Hvnf6U2evxM6+aZLGym4fFsjYPeAr1Pl3TaR2Q2Ol+LccZ+pHLOSzgTFaqmYMQI92
KnQLSxY0Mu3Q5600+KsvSO5p27SdW8CJP4sZYHGoDywSSNMKHBgpirwjhayEW5Plb311D+ZZXEIR
a2xpl4YkKEZMgUr4QIWd/MEzHLFUupmzR7yAmtI/pFkQVWcvJ8wFzf4Nvf+DqH2pqWoXxUJTlL0J
E4JSGfSmvk4CX0VMSPr/GRM4ZZAdE0TnLNECKRMW64RNnszKgWM4tbHuPKFKjSm3Murl4LX+BzsR
wshDyGVnxkOaJtcHnMBnjqYszsQPia0T8Umsmn7wcsFtcf50f+agnyJeuUd4ASMk74QYc0ikcjti
lAw9lu3b3QtEt6zf+DBjTvr/JvRJCyODfRN0wh79T1ezy9Iqjl+slifV4r1frGb9O7zW+c9FVnw+
W32PmIlt4uIIBNq56K6BqmyV249X6rXE7K+yI9ozDCYvPPsYwOk/SYLEUixj7ALMKbZf2dlqYNfa
Au+Z1SPudoLZmpUpN8teqq+lLW7pdCVC61ATHYKCP0m8KOy1m01Js5+BvapPDiFzp8KeYt9T2e9n
OCQ9HpwnD+4xinOFRMthICjHrEJEPPJ49MVn08tpOZflzof7LsJTJKo5vWCeaaCZVQcVapX8kmW9
ES/KBDEKHoWhjnRZmIqzr+OJDn3eW81QX4IZ0qIVWqyOjWM2Y7wF1r2aWe83dLPW7FrxiddaBEIS
FXrKkeH3zX6GkSnXvhAPsjWdrRf5Tdu8Du2zG17SZeSsJeVdyF7vkJhOG4pO9tvax+6cRa9qQ1Of
tw4KEFpynigpvBL9zmMO4Y3/RXQ/Lv2ifGnEe1b03vqmkYukwFFgVsBOF33qSia2TluFb5+p1cdf
5iGkoOZLLBNvUG+PJn1qKcNpcahXPi3So+meGOGgc880aIXogxwGQK/XmdoSJjsUibDrFc1qxrfv
MP5c7pwLMT0ujey163/SVpPpr3hAkWadmV8N/rKlnHMiAio0rBKFBa6dr40pnodEwresLYXbxmGP
8pBC/Vu3CqKlIajvRWGyIbF9TUHpenhc8zWfAS4D708j2Rdanq16o2DVfWV2gWZqmVieSbMKCzDP
Az4tRstrx2XFYYqvwuDOjF6hlcmTaRqOlgxjyJOzxXBR9aGBaXyIIebcdORNfRqtOrC6IW6tmJP0
i927YolUNfNpQ4LsYT+lrRDdlHIqcysavTrf8+mtryXl9uNwu4RofqslPMmZBBXwnXYjrFS0FMh8
n/noAchTgwDyUSDpuJ7OXHplucyOAUyppurUb8rP0dy72XZQ28L8eMSTJRZzNc6bul0Zfopy/Drm
Omf6NKToTHeJ+1YxQTJltA6Yhyrs3CIQL9xWlg+PFbh1fnXfRMbwuM8FOpkylTNf5t6aBXYCIwCQ
vuMwIVkJOOjsj496OetD75q7gQjIxHf8TvohLvEUMMOLF90YkKJib5L2GB9778Vjw6B77mmjYD7M
D2SP2yKorDgdivl90VMeU8yf0aQhIGyIfyi5oI752l5L0leKPSZ8+Ym5cRbAjFxsviVIKDvurG5I
VVV0speLTlfk8aN6MLmWKJTWom5MC8OP8YC9XXx9YinRoCLdHcF5xNY5IL8t8JUrLnavrZxTHOcP
/LfP4mEejAQD+tGtBcy3mSZY9yGyDmYdiZ0rp9K8KkHW7KkmF8AH55PidVe+/J6W4oIZkqlYPWy/
XjjsFSKjKyWuKdlxKuvddo9yvfHjCYJo9hIbbDYdmhIO81BnrLTZwgqi3FY8HuPb9eU5cVMxLeza
rm5ZTJ8efDXc2/oJhGrc29Noli9Ggb5iSYq95vDN5ZjlCJo7Zn6L5Puvhi173T26W0/1QvLhLwLT
k7IYnwMx/3DO6ZEv+T4tOVfy/XlM63SHN+bXAB03cEJYGw2HubE3xhvJd1fI5ntNs6k4bHKKSycT
5SIsiumo/p7ahBwvfj4HlHvPu9G6xtxXRvf81JRFTZHNrbgpYaBdLDwl7fALxqUixL26tuH4yMdM
mstNSGtkI3HBgcx1RbbC+aPsvxdoHHUwENI9raIh2/KOACuTAoZ142wY4/BMXf5S370h2QPpjBrr
D1wToaJGjMXdkbkQ2PDGRnhTg9IMJ3NMeTt3VlcWI/kr7LgjTAd+T/cZCsCnCFvkkkWhfel7fHHN
ridmUxCIuzpybMj2Eq+10aJzjH/bFjI6B8mr9UJYsNSJT4fAP5vl4SH5nSYmmq73c9I1mCUysUd6
W9lvXyFQYcCPNSPOVbpOwZVklrytq1r0F3uWPeVNUy4lgEQ67CQeERBADgn0wQqvrXV3o8QcZLEJ
LjTi+j4SEFx0kvRQwpGLug5t5CCYsQoV2ZqQd0gOIxNOKd4s4Vodes8aAs1S65dukuNUTsdVajvJ
BybeOiviNed0b8f3ihbFckY5TpRC5cEFIAF+uR/N1Rdx00DWGROBc9ZO0Ly0bEAFIMJcLR9Up5FR
4WL4mAPbl9L0zI3f54vz6dTUQUj4xUu3hRouZVgWVlSTBmEfpWuCnjlAWDNe6XZz64vxWN0xKNME
viI6kNkKvs2f9u2SACtv6IMjKbQPnJmx60PyQ0SGVsE//GhEIByqbuUGe7UGO5UYpQLCjm+4TGtI
7hDCTRjxdr22xL7r7ey7tMbsrcetEH8lQdUmUR+mu7uBbBodGZVC8CTUllEcXjVw7Ybn82z1rKwD
J55sc3G52qR5QQkj8rABzcYGVHSeCXUMgNZRi5af1N6HgdEoAcKqkuDeqG9bOCq8E43XJQULvcgO
Q1mkVLW54sF2Qha1r4494KY2mo6AydDBBZOp0qMNu/RL962dpfd317dA/krkZRaGZg5igtwfN6Ia
2V38/RiuhhkEsh64MCw2XpfU2M20t3uke4kaKmd4Xj3gP7mOulBtYUfuT/FGbTGgVUWe2Z31Yxs9
nLXazKE51spsWq4Qf0Ced1hN3d8dGIZB0GNKMJBJgKwX9Z+apgCi+iwPU16HVYOfI7i8wY7dJv5h
OVdtC+rI2h5SAy8A4Fh5MkicG5/2KLRC7UQxZ9ynfcPqTEpSdCfhGByk+oKYLD3bXB0TrVV3KgCC
nlimY4BOnYRGsbnMGYkt4kL5G/kb/AnJNW/4pgHfOWMFIsmMF77sxLLmaQXwCpZodaDd7uGcBuwz
RTFZONKKxPGsx2IMPFWT7j67ngw5f5pKQMdLiy+mSJjy9yfg3zDhaS85wQLeZBQTK1qNyBAqBvLs
u9qjS/iPn/i4z+KgRfKa2i3p9Q1n21XvWOPEqdcCr38kjBl5XMRK5cdVi0nDoZpLa2A53g02B5m5
p47MlTEzLC6Tv826ctcnqUWTdUehIHu0eJr6QhKMCoJ+AWMx96FS6QJ9DfY3Aj9k+HACsU7eaMAr
6tXLgxCLKGVOdthdcfnn052P+Ln2QyK9mLpArz72JRNdrIA0tZaZnNCD7Dbx51QM5Q+I8J7dCrnI
fZWFA4dxdhumaPhW7o0m1OJX3kxX79zUpQg2sysy5Y1jLUG6BcWm58XXdYjYR0PbFDBh5+qrULmw
IP+pM3Ee6DiR3/PynGXBFlgRazAZgrc8mlVTbUGcnmTxBf3IGd6IcARpfj84pISFVQ8mLZz+Zk7x
vrRazVuWDkWCyuMTjXbjQgjGH2AwxMmNryx9q1x+iB8YUErV1JLhPczHZbBl/NylRHfd7kRCFkBB
WVfapBYNZX1uIwnHyPZ8kIaGRZ8W9ZG9+C+uz8JN65G3XSPkSeiMdS8ofa6Me/WB3nlgVWZklKwC
pUYCaz6VLy8wOCsf5HId5KJDRZC1MmzYuHjtwvHPf9GmuKKUIMvIbFN9BQyjBzdERGShiYBlgXME
/1q5KBELiku+3aST0dCBv5gi1+k/XY7yPIxeLgse4aYWWkMkrc54AD6GzluT/VpFH4Y0GcIYybDm
zsxl7fiG1+eNSWr4f+NAd87ReRcVgljZ/8r08lYz8IU0Z7qQm/6bFH7DFHPB1QuHBGPtV/tAjiou
zZPcTLBTSzUXj14txTNE8VJ73BoNO28X8qS0MkYTIzAOaAK67UyPfMUQwoTubQDu7E6BptfmZy+m
zhPHAxKYno+63ILwl78ZP1dS6yqs2VTrI4Yik1VXA2oNUInoq72n4HQqtS581bz2l9ozgDkBck+x
j+YakEes6ikbLAQWTgRebh0kH8YCWT7taavQd2zWs0EHXfp2Zlm6cVl0GRxC0WfFEi4XgWnt5y4V
p709ovj90tm5pJUnLwOPEpyaTwOIl0R8bkYdFQNi8yGzs6TuRB69SaqYdET+UQGEXTedFBWjSiwj
bPMXZxMxz34a1Ar6VvtB3KWwyXGcxuW0tpvrE2rAkWiH80eAi4fqf2pKJpEr+pqyaJYkE43viJRs
czYTLrmSa9yKM4W7BKCPtv+DsqOxKL2LSTssYWcYngtc2kR5kAR3tKUJCi4a/IqkmpU9Xb40h6bB
0uLdEHn+vwgR2k5ZQZxfmTBGT/51F+fUdo9nYVySToXuprDQa40dw6QfuSQN7a1ZK586jpv+Wa3F
XPivFyCflGqN5tPK1GuC/sjgu8rpV51FeA+NFmZX+0lMFTJxHdwy7N8yvWpUnUCaaCKEUS3i/RU/
61wMavQJDaTByEGNciqAboU20T7tmOprlT/JGH7vh7jY7oFttDY5JAiaD+0SX9hun0+l0nuwbgzA
xVxtEAo87vboxkT2TjTLpA4tLs+De9etzREqkzMhoMDBSKBLIGj58f7WnBFAN1Tw9k6atKZrndma
iAhgLxEerDOygNGfHIvYisa57o6rVdDuXJQDFYdcSI7VJDhvINvK4U9xPebH037TJKURC4EKjKS6
Ij5eRAoFZ/gzMYG0M8bJ6PBWvu18hVJNgAui58JurajUgTRkpqV3SBXQsM72c9/jAYvTEFp9KcVS
NeMeo0vsBManpcQcaphw6voCzPE1V6p0i7LcFkgw94UtbY9Pe/DJDW037BPlEuc+eipp6nuqKTYY
KaPrq+0w2uzPf+2zKcPKQpLbMxZSkkr0QH+i6BfFLywRDu+vkydCQP9P0MRY8z/23oq7JlH4jCeL
bYskhuGrvIdSVivYxZww42LoL8z4dAFEOJ0wVX2gKQUWb+X3pu52ta0bqwyRnJSGoQFrB2xl+VDn
p64wf0QbvoWQ3wGLkQE0kFLtpg0JmVWZ7lIN9mfokMYCDF+MgvAvzP+NVnva2aVGJFshC1rJgx1d
VHgsk9KF+NX94qZ3rpXVY/yndEm/hKGQ9aKgrh6s553TM0AetyEeM4Gh1qGzNnMNtGRoeuzf2q2L
86EAmgU3mYn5/7RD5FxoGXmXP+kw0lERygbDB4ZJLYRiX+hY6hbFSUAINV9+sUY6gIRme73qyeKu
wMnTguKhvzKOSF3vWPfQAyHV0IQRxBqKnsBSxVwn+nHjLKqy8ijLw1OATizOg71L9mmx1MqIhkN3
/nhP+RoWTkvWT31eCUx1gtR0xWe59z1fRTGh66jgv85aUWVKpbrpqJA/K83wgb3onP766DZrlHwM
B1WLJXSUO7gNokda+ytPEaoTBN0LIQSmGx7hUPI15JKXADB1FGJ9hsqpAY1UabtsIjGTVHCy3/qP
ycKHKV19A5VtSp/K3b6DbY0qiV+6owuyVN0y4wMJtsyrFGXP10LlO0FfpJ+Xo1safaHScJRLLJXs
ixB4j/caHWc5C/ZN0ZDGCKS56y7fJm3lekcJnp1PvfNvFJzXopdogWfk24Ls91tJx7U27AdkWgve
K2RdLuInU4aoTlkeHOpSTogI+53OjaMVi5dFI3uk3DUi2Kex5TF1SsNDjSwkTymxbKhn4OGk1cMy
FDIWWVNhsC7JQc7b9OemQXlFHI1VVtn99d0fZl21h0F4svV+AQkIZx3HGIXsFLCsFXvTJF1f9kzN
QzhUaeQaPv8ZRVT/CKZpB5s1xGn0I6hrTBTvk5TUDjrI8jtevlgrv+hLk0BMwBl/jDnRCdX6G5VA
aUH+IQU1MCZk1WAgEjG1YJxXSS8Lcyxt3bfvl4ih4VuFM6AgxUEBYbeuIVVOgkTxY7bJAHvKQgPs
y4LTnQQlA+eBPyjiCaeu0JlY8ZKPpiutRA3ESZCNSm+MD/3pUJGfwLUZeR4dyFYW64vVt3NrF0BS
57ivYjo3c90Po/elkt5gnbE/GI7MOZZQpeqQ3nzu5kEuMsQdIvsonHBWxbYD0ZzldO1GOg8OD50S
MQAMPLMlM97/nwihreE7BboB4LpQMWbsM7iXSEjKkikL+QZ1X8wKLa+pwR/j/l9sDX30xIpn7ija
mspqHLU/TAQEBovcC08tsvB9bvkczCCW6vqSeSgCX4TRZ9PjVctZRk4iIZWoKgsynH2znb0KigzN
wYdwSNP0X/UyF6ImP19dvbDtPhkOi0cDoKWxBA806AYIq+y1gccdye7dUgENiWJwUW3dAxP8xggy
QlsquLZmIMBBJ4OkqHdZnyZHC+egvfYhWia83CdHbKKE2Bke8GXgroYLT/rzPDhOf1/y4DskMvQJ
JRH52tqll5oNXYCPbZL+CLAlnVxooRITPrMiVuNH7zAK/Gf/rFzwzTYgbKlQ5108yqsYbWLH5BbQ
YkT0bMqZ6h6tdp0oUHETd95FssK7DuBnlLL4x3j7+F3VUzd5PilqHoDrBugc7d1/9Tnre2MVWd83
R6qKhfkPBH2Cqod1WW9P0r9UGS/cpfPcP5FlCiOdA/0HbJphgW91nr6LTxtbPfmP6rdJfL8218F+
mn3nM8Mj0ZUBc/G3x6ivyQZKjNnu/VbY64MhjQoC4zt2U3mu6Ds16tHz3/NV3seOqmW07K0PQQgD
wxB22m1dQFCL87eWKdAkgMmz3cTtN0G1n3wisaECKFSmN6tWZh3f5xxpkFmLrV+0OppJc/yEIoZu
8fseRv2NZzaGgH/YoXKqCC1/lDwHwp/+BugePxA6kTQ+PFktAiQhOU0hscFnKpn6L6GjhGFbqy4E
4GRHMyLwMUrI2U+iAGl8lah4ZjEB9xKLb+8IaQSFWdiXSMRe28Of89V5Ejl8SD41KBKmb6mD+l9f
Ixs32fSiuQxIAZ8N1aM1HFlWRECYcjZitcoeyaGomsxZf+J7L0KnBZ4b6MpZpQToR6DavebKO8gj
UzUtqGjX+hwgjFwbm7r7H5gh8lVESDfl3k5sxS9Hg2Alej/afuhlIGGCZ1EtydyuwZWU66DH3y/T
ITCo4undiirfiWtm2XlOzAJ4jeHfU+EtnstovfZKlW0Z3WpjhD/aG+4JulnAmX4mwlRxTa6Tq8GS
trorGad223+12HdBN9i/Emmj6s48v1Fa70uF1TZdXB+qpPUWFNmx5Mi5DY1nf1p1WufEXcnxDKvG
rcSwM1/YW4cTTA8qRGaPVi9rDaI8l5qrppZf6myhuqGpYRnJCm0+xGv9/IspIwlzmOL1J58vo5fS
2VJN0yM/V0cdjueZ+K+nwXAAwimewIZeIDf4YAW+o7RKDhBsuwfwV2A3vswcNJY/MgwpoBkUBo73
A8uzajgkhBslmwGGSH6UbGeZhHHun3amupc3zSecAG03D2clf746Ga9/emvZ8C2wmZYnhDwfeMW5
JXzTlgZ/umGvczBWtnqFlhKpStiPp3YlWfztHyg3qUNLqnvlzMp8/IHpoTCYyZ12veSwi7QdFzh+
dPSb1CrMNrHBhOzPjiC7FONKqxRGeNxlOFXqpWjFTekCmCi4BQ6375hy81p+GPvgRd4F73DOqjvM
ebAeSm/oWCqIzTnICSum3MBAx6OUWx+s9PESMMH89NEX+xHdjMYmt7j7cWMRdf8yeAn0sntpGDK6
J5UXkU5adk75PzJxZ0rcQw48ehzWzdMjE0x6BlCiX3EP19FV7b5PHBtE9X5WJ8lsYujtd+M3zoZA
O2EC3QQ5cFJc5umg7OjW6fK8qMHLzLZj48siYEXesjrjB1TSa89U5ZgDkSzXAgCdNAYvNwSvST8J
7ROUselqlzpkcUCEj/dgJFOrqdyEjlp/lhpJajyUVozoSMo8miiB433XjB7lzR2AXOvhtYNjxchk
lIqpWUJ53uOoKbn5jIHzC0zjR1NVLtQmnapYgKXSth6PiXqKb2Tug0KIHlJtZvQda4QIsHe+FaQL
smiWmP8LjYHxePJ1N7+BFWoWmpoLvvfRFTkcMqq7zjcqzfY40mifnqSPWWTd0IwPFtzq/5oSad8K
CsJ8dfEsSb/+JpR8GjzLF+7NP/VFx+l8jrXKF1RsVhV5Pw1CKBEWP60YIXKCz2OSYyuCbpVzXw/G
z1tl0AU7a6DYjn9sTsij+xpZTOq9dffDgOD5byT+BwfyUfykoTvMFNfSF/KnH0KOCdpuKMx3hnmj
wT4AwLdFvFFFzmO2mw/1OCEwXu7ZUC5OqibZC0sd/lmm9qRvt8CudzFDiVLkyZTrRM0zmHOeUDCM
EPTKYk3qXp81euHSi5o+0HXpRmhHi3c0FtslYCnKzvZcWQKH82vimxa96YLPoxSs62sEnKwfDMk3
244eKln2wzWWolqW+mPvzts+cLXgzM2Ggp3ZzhbTOfA/oPUa2zV4nhDnpShW298NvQoEz30LB35x
f7CXDp7FBouHNH4p+rQvkWHCc6f0TT7HcyKfnwJZtcF95WpYmcjJp/e4qJ6V6+Raz7Fd6ExVpyUO
7DwEFpY/AVpP/1XVgl0TJTn9//w6sFkD6726ytlpPDVgKSwRF9in8HyO0HaxPskCj+/HC6lbpj7L
jqVWBmZH24f5W1l2IVauc26a2UNO4oy5I0lH2NDXxXPko1UoPii+3gMW6YZjuoi26wNt1EJiNPum
+oKrmGlD/o7QubajSVNBKvRGWiAkACevZCbsBT39mSDnhVS73iqc9JY+Ty9hpiodexXbKLA+0vPv
ouyZaNo0UkxfoWW6bvzqg4fisM20khTlgAxaGXl/TUIZig/VvjSGYbGH+qR+IrPPHoJoBUUw0mxE
lQ/agGYwve6wpqAp4/3GIA08OmVpOjG3LC8zCmDQuFHVzCH5xBWSndyRcs/fi3+naHtxY2saAwPX
6zS2dyoKpVwYaBYx4E6upIIxoL37hFwBLmRnoO8jA82tUmfpx/aNxnaYh89/0lA63SGfwvlzlq6/
QY5GNRD0Cwz+7Mt9HU8jzqdZRFvyepx4Th6jBhmZw3gOLhfSDldhF4G37ONkE7QgqNOVIfLOMzA4
3Av1of4D98xXfp8+5AgXGMotU26+avfnjmIIE3C6EDJ4IdUIlve1m5m0tsNN7usjgmnGb5VgyTjA
2YcAaARGvyag/7TWN0+/ga9Gs4NPv+KvQvMQf5AlMXKTH/abrh+YVZb2lrsSXZ6YVTOYnZVxiqaV
a0phKlmWWR3UoAyMxkJXEXfV2eormH0+6sPcxp+KZQxJrew/hZZcQ7NlIP3i0H2a2HcSC9y13g2b
VXX5az6J9nbc+46ksTzANfjYxbNuEyUnUtEC0YIsQHkzQG18KonKcweUWM/y2ENEttTXw6VMih3X
7e3B9L3UVa9aJd1sVtTCtxFOM7/b94Uquc0h+3Ckm362L+rsveHTmjUyxHD3qW/wchGiZ0OdzDRi
rnrntcRz2X65MzTyRHhb2dnw2P6ZkHhjzxfwCfgDK3nfV/aXNswVu0ErZ154YBhUEdkU38b3r1dG
BligjJcCXvZMXhG43GHUK142ElLWg+ETklGaMzUwBa/5zRkDmKPjjatb89NXsW7WGPFTtbEKq2y8
VBrBTnIPPreYOMDiHVxRYCxNx9Yido0cPrcU5rlzQME5YF19aq4Y/RGgN9z0BvGeXlEbNg3qJ60M
kmJ3D7LEy4565NK2UpEaWc+GKc/wZvlN3ILVL3VnUspXltMMycGZCmKrM1nJHU7x7YGeXCokhg8+
onw8J/1B3xDWpE/2dQjvo2Foi5nmWadquApKIzbHrs/dYl8NtaR8G5eQEN6XD3piIRZkk+02RqsR
HqiK7ZzGwFBNVo93Sgtzcn5jzSRtH47cttp7XzUGYnOVwHwxKY0rd6XThp9he06FjzyXTlrDTKgj
8pJ0em6qB8/f9T6U4lTu5fJFugQiYwfkovd5D766WO8z0WYSWLJQfkI/2DXNAYRAccioCuINoU+r
/LifSjDitNAkXrdUETvbSioPZ7K4bQD/WLHUDVtkBdiPGAual+cdHZn7IAYqqE2DZlrMZv4661Ws
1sTEZhH1L0OJB6J0QKLdeM5Ze2dnl2RNMyfKmeKL/jgv0V1qHj4le40pf118ieA5PfXmAMMRleJ5
U88QkHdt+I965id+1VM+eYk87x8dS2ff8B09XtsZnut0g757Gsd82TOgzlFIestc8pezSNUoIELN
EwObilLr8l4LuZ+sfGhGkXLZT2D3mLbATchh6pa/+6P7DE/xe/nJhqvmfmXklL365G24cIj5UVV9
kiVhCyYC+tYPca3H7TlPmG3hAwLGcNBrBXOCONE6fhJ3tv2DjltwIOEMOsCSZXw7AS7QgfMzyxxG
vXger475r0Qg6MS8AqusrzR4ppe1UhZT6qff7U9Wcn9jWWBpLU0IyYLJnSVepaEEZQ4q6JbxBLH7
Ct/xh5eGanGL032qmQy3OtUcIGp0mLY6wYWGEWh5OWA22jZLtoxthhPQMjfWB7W69rAi6XOrYjn1
inP9SxkfS6WH0w7oODpy0JAWwlyPsvVIWJEOHc9VgAJSIq0YlUVRX4LHD9ti/fY+X40QXJ78jx3n
ISNkHEd+o9H0ds5KEgp+3DlWiCvm8RQvp62Nu3tQb86G3pOQoCyC+g7Sh6nKvJTuIHTYvKfcCgiF
23jldml0irvBU9ubxcA6pSba9eKyZATg6Zzzzp9b00dkzyiKY1KK9LH0Y1o+QbsA/pPk8rSJDy6w
0WaQz+bH28jBPdek2fCA7S7W36X952hcaXqRSvf1ltcDrF8aAQ1VVvK2j3FqxLWzp3jSAuds+BsZ
v2uRyBy2MdZh0KEd9/+AGqFczxgsr6rnICtWc1dO2Z54SREA29AyyDkVSU4SNDRXvGK+643r/6M8
JAOCDFlnh7xSfGzwBbSy+WPW0/cMxD1zqHaNB3MyUwSZDP8xYnbRYGFRx5RxFDXIpYGCFfjTIUwD
Sta7LixwkBLxSMT/fm/UJ+vIaoX61pdBJBX6x4VDVOQELMMZ3uobiZYsJm3cNb6y9sgO66YF7o3+
qvxdGg/DYKrbPDRKCsnwShQGZ96SafplT2CTDHSVbNmEDWJP9DokaBtzgZ9dYJFZlYVAtwACB6CX
SODNGCK489vEJJFpxFlyqufrrxcJwz66G1UUG7llahvvU58Jow5d82R/PZ1B8GzV8zSaJ21/IBsx
zbCgnAzgWRWFSXMzBvKneDSOHbFhrv87vbfu0yfwBB+GM7SyVjoPVAPRkQ2T8MxOMs0t/Vk7TuBx
UcrYfhrYhwGHC+xuW0QYGcTfl5kVmq0IR0QjgPxVDJi5xUrnLq6jjQMsrPxulptCsUw6OtWCYmUr
8EWt7q7idzylvaw8mXxB+RsE1YmF5K8PKSc2EqWDykB9SAp+wA7JxZGOu3Zs4lYsC6heVsvn/g6C
2ym1TuIftX+tZIHuS7LHNKSZ3bH7IccqUVi0F2MvjlRNOeRxmNnqN7VTeT1KHE7V6Yolq7PsfMDy
DrAvEAqJMFVoo/3nBAktUJanWt44oTV5vdhXww1S4RDAlKsmXT2MVT7/buZSDgy7gTWdSWO/NRZL
PRRJ4zxILisvgtF/ZCqeWnNhE2E3zpw90Ccy+Vu29CxPIs+IwmTrBS++bEQC/hDzoRcaKzp5tC+G
Zdss8k/E8qUD8/Q1EfSgzOaY8N8xwORKdBtZBjvKi5JA2zVVdRmstj8/RqJXbNNrl3I7RLH/J7TU
wydKM3bU7BUpNETFjBi/nyRBPzIywmugiqxcvcuDidnWVWqIMilHrXIZLs9LkN+DRM/FzWQKZZmL
8817h5LznMjJ06F+n7fz2Enhlp/X2N8tIAFRFt5jJ2sfpgSRyV+mzQqNRLT0hRqlfuiG1ehhphc5
doxPRegjJFEehMzOg2cnszAqQVuVunjuHcpQw7RnSPvqhBXk+RG6FIymFeOnuKtFtkarXc9pqZ9P
qmHTHZtJ6aMkyfM9AL/RTgL0zhbDZPBiBAzxRcMNOSXAA5bnLV7RdY8WWIbgDHYZAiZMNw2V37LM
LiouMlxi05NvZ+5NnUHWHbdDNJb0aozO8Cd+v/bC+JlDHeJnYVro4kN0WeeHg5gGTFA0JWVLAE+y
jiJByohv5uTBgJXPolf0Zi6gOWMyIKWwYbNPTk8Hlj7arUM+JU+rgwMl0KYXbnIeZ9xiBOFnEaFN
dv7Nh2eHfpf1n0vo/foNE0blOy3favPobxOZDoikSOaNYMeMXhjSFzWp/SDvDokzBDiUrd63G3kK
cNtrSai7irYfSIP3CK/jkL69WEe/hmrNoatu584Pw3ShUsrO0OxK/FoR7C5tg/9O3U24t9yEkUJx
VVd84ZzGma2CAUuiYs8em9z+6T4aJq2qUBUSXQyGZbxkUAir5opSHB1Kv7NQTlBGgZXoYl9Opxy3
8k4PwaDnce/xeW/iFkyq36NJVLe+3MvY2L+xx9gCCxcecxOjMxGBYouSJ8LZ44oCvEz4uJp5U/BM
hWLJOv0TTHSfL2EKuqu6an03h4K+pzvUyV+Rfdqt9whH2VYcJlwPRC8mVcaKyZFRG0TKp+oomG+3
C+vvfuF3oXNGNR9M/W3gi2xlfrMnJfTVKG2WkLOZU4Tcu0kTwLfViW3QhOQS4fHeZU+fX1utTiki
OcFhuP0N8JBC7xH8rqcA6VVXHwP820+9wnOoNjA4NY/6y6IgiSTJkogC2nGZEB3kmZne7Ltehc5Q
IlTpb4aihVsxzv9gQWeTT2k9CT03aKeMVWdcW6ET8bhI03Nq+26VUAGKMGL+DtqAFIW192ctIEGT
EA3bkZwFoWtK7ENk9gnvSxJwwlCpmTdSqjcpHoz0x/K4SSMVOBjr6xj86zJCA8ReJYQL4qCUELlT
6/H86jqwrv1AIMLdNjvoC61PGnFah3aVx9NQN/YARaqk3ZqdPnzJQdoysAfiV+ijnlN6Mwt6j5Q7
qeSkSrBMzCDt4OhWbsEQnL6HJkzbC7809XlBBcn8s5b4jtKL1r4mJI6qbg8CxEbcMEF+Sqpz7pFm
0t3kYXmJH6NY3txuyR+aik39phbnzkEj66McQsHOiSlMxdJlx7sEnW45WPQ1NUBTB1unH6jqdppa
5/QQjfAgRjz6Q+XuQ04eDuIbXn0Bxj+XLkkw6zRbiCyFiwoyyiDakqQgbegP3wjAIBSGFmDme/rY
L5/eupftQ+rVaIxlNnbAarfHCjBcPF8CfKh/78+1Pla4ffaDkyZPNoJ2IL6hzqrWrREPgO/0Cqke
9CYrfPBFYH+oefU9Ii6kWpWTyGcPnS4Z3uJiG1v20cjVv0FFbFHGn3N/ltoRPGTfvBbHuU4B06Ew
GNi4wf0ROSKZ/q3G4HM9tnddApfFtEQTE4m901iyuJJfuKCdwoSd19K8Q8VXTncx9Dn9OPuhacKu
suKL1JIjp3y5FkP/W2mh+As+pfuO3plNb+61KDI6EFFAzDTA3DX0TBCwApAUxFKAFB4N6h4Ts9zc
B4uy9vm71KKyMUZNT/Gl3WMbv6PL5LYFsurjuUYt/tKQ4tcIopEzXPA2yyIiBMAa/RR0oxKoJ3sn
+UN190cQo3OYnBBkA0xSkCjUhr2VX4BgCnI8oDRWTH0YDQzIPfazh5vojqK6FetSgqa0+bcttsk/
D1osXGh5xxndSmeJ27v7x1VcfHo3n5wvYluAIEr5qhb0VJfEsWXbLVBKsfYrzh+qIx0oe51r03VO
Lca5RqL4qHDnIW2sgpTxb4KXozw+Rb0Vl3PkBo0c6ogqsoXve0NoD+t4RkR+f/RMIqRxavqIgnnH
CmTtM6OduMwtqVi73dJMUnWSWut5ZQiHvPFKuvYaif2oxKi47P7AvLzlwTew6+O6ocaRKlva2TTW
sIfnEeXHJGBTOvi+Qk3JS4NQ8Q2TMSAVgvfv8ytyFRhf5CnJ+VfPvthCLGoaDKIqhswDLc2Wydhx
1+67ZMskSb8cnXb6kYC9PsCuDbC+6pjkRQKJ4kGHhRnqRLPpTTcTMrnsWr6WeH4FZJE9fcSO+8AV
8jdFehb+hvbmmYMLR3nzm4kcunXPpa0kT91GufBvy1ybNCzmvFRPtprkqo9z0Ts0uxOUjQATb2jE
CoWzg+nahE6HQYkjMbV7gy9Jyo13A03zR/jFXAj07H3MDW0T0MJoDRpckzH1vMijIwafAtw9NIbz
efjs14vt31dc4iFFaIichUzcvJJcLQuYivDD1L4w6tpf4t0F08ZAUCBsq9bW/DblhgIcz49qwizk
Aa460yOMBD/kbbjczYPxDvV06ahsjM2f6wPP44jqMji7f9RBkK1kGHqNEYHwV6SvvRChfAR4JG+K
Dpo0PASxjanq4piKcLhBtgl/bCli+1L1f4X8AFlYB0LZ7jVhgE7KHjU4aInm00KCnGD4nIFlLAIu
s68GrKBTnTeC1gEMBZwhLdymN9l8US4o4cfzxLR7tpSum/WHEtbPqNY+xM6fTESo+onNl4qOgltR
r9hFdY9DEj4L3U2iof5FbmRRBOS45jeiEEKlr03EwzBg+XZmvpW6WL8R8ipSriKtEo8nq92CdKY6
NTz9VaacnCRoLc5mPn6Crm18hjURexnan8lLbPcczZ5BrknwA6eTia1ydQAQRigAhdD2BInXXElj
hCaJHsgiEU+8xc16TZmc4GEST2PysWpBzdU7EhPggjxgRdgfqWTuAtQAUIEIv1Hd6jnGrYqPlSVd
QrPHSxjtHywzUPKBN2FN+1G5Bg3/XPyU3E2dmsG4GDkDy7lGDUWmFWO2zLoL5eFTZcGBy9zZ1Wef
rnD9DeYYTsOI3tddKno3Vqg6jMWpP8Sbr/WG/4tWpRtdaJINvuSe/qteBRK9VN/VZ7o4Ba2TLeGZ
3w+rvsLX+pnBi5XHlaSfZfYElARj5414tBtUO9p5l5CV3R/uCrA315KRe3X7HpJJxwYTflS5BogS
qMRfJ7yZ1KOqJp0Uv6ZXBANmWVWCMgwbfl3PY93UzjTWBQWzxaZb7fqCAdByr6O3gXOXMSCJ8Oj2
xaUbjCwwftuMEfWdj4T4mH8n+UdCU7VPDieApD1NEtC2kCvtEN+UEDAQEuOGW1dXz8LJ2Og2oX64
hDmWMnmokGAWEXCCUE7cxf4KCV91RZQT9Fe0nJ6oJDM25/agea7mjCEUspNHTK0Udsnc3UfVMXT/
Xr1WyuhgnRp78jyRxQLH1EkCnJLmjGDIEnmypD+/C8y9bn7746hZggFHvnrpN6nEjXbCKbEjYKMc
hS27rYj51gAr330qOiCTcs+M5V+uOBm8jlcliL5t4ThoABZH75oCpCBg0x0P3/IVKhrHHRzutlWj
lzM7f2mzdpexSqfj4TpuExZAwS/YIgCuvy7ivZrv6pCXGn+HtI+B7OLOVtJSxtP+Is2XqhCNC95I
op4nBCc+ooYGo+CNZuukct1+PBuyh+6y+TWGoDmnfBpaeUPbGcwuD6hENahiMA7FLBScES9YM8rU
pEQlnAseORJekrNQFWmqcwB6BeKXit9dmPpsViAMF0h/u4gQlTo07833QFyrJKciGH0qAZl/6WbB
Nwfk6RQp0kmPaKonFfq7QqyGwoxAJVWEVenkUXfG9qVWa8ycONo87IBJQhraKUW5gQmhKjfTfp81
zoKCVowJpefwwWAQCJH7uvBCfhzLuRlWI6ndqVZ8fawu9EH+WYpDdtL8Vu5nk8yEDf5I22dRps0F
9TX9LTQ5KLoPoaU8VFTmamQVDWYPvASd3dYAo8yrezzUMjE9gMKzBGUfbhmEjSWVF9qVay5mbm7G
Pa5JnUW/6jiC2ttxM8R/XCskZu/2K6OcOprBytOude5/awAtZmebuDFt/QVySz7x0FZAoEjNVQHJ
D/NjgDELnEUUsKkKDs1gseO+ZYPuJsalKFUohEDeERn2gz4Vfih/TvMcdMrsf5PNGpFS4Si01lf9
DEcEnxvFn1GK7+Cs+b/r+/acuOR9b0APkPV4dbVhp3+UrbBd25MEDxmwvEaI7zwZHR8BSuDNF7+G
btJe/8HWJ3Bv8oAGzvVtSvRltX+lZqiO3ziho9duVuz5Uo8VsnaHB7p4iZxJRCY5dUnHW3BRY5nQ
Wc6qcF7yMXfnfS3OnLcgPxkZRurjVaIDysI2o0S7rNPXqkq2IPa7BWXK+0Dn6phfDqrdkhp573ay
WW45qvsQH45c3idPinD5gr+S+M0p0TYjywdlC6n2X5tPFuIzb/Ocy9uOHtdlZX4LLecol9cOdrdZ
W/WnuciGgTjuskCNCR7nXccARJfcBEYUpyqiZni3UeM3nQHbxxMe/1PGy0Qvkw2jpj0LkWspu1f7
74icgMn9BII5T66mdzVVGMEf4OzWdp8umZ1sRdtOLf5B/OyQyMpGafreXGfjYHiPhfRnue7C72aN
gH7+G/uilwQFwbQJzsr+VYIpPB0SPKw0TkAAd2u4jof6W/G8FEHU8EnKGUOHzHniisaiXHTspqln
HgV5vdXD6M/pV/2LAtKFyn5Nie74hyfhD7M2n8bC6zF80uAwqnnOA0k7A7jmGamK1/zEevcddC00
bW+Xx6aT0r8ZNOIpnu1FMaOAWByYd93tJFrGjw7uPR8PIKK1t8p6kbbDkQpijiMlS844akIadwnF
Oy+Dn+6xBa7xTqu9X7QOt21ASZqT9AT6+dNuFWaBdMaUWS98NzyNE0IQ/a91FIJUdKfdpXlc7F8W
oHUrwbmTDLQ7R6xpwBA3tiHc0K/qMmkNRXdOwbsI879NMMxqGtJl/AZ3okA5sIVKgqMxtQ3sb651
gp44UpcBc2ia+453/M8hBRVD2n5n3r3d+GwvBuZkkeBU2u0G8i85ZbHTulQS9J7glKk24XmzFzov
vPJwZHA+oetOoR2uDVL7cwNnFeUcz6zfrQyULpLXIqZt5qyJXJ5PTGwHGVHiURhE76tKcBjhB4zB
hc4tViFrTXk2f3o8XMEIqzt/eUy3NArldoUNn9pWnODP7YWeeTHbG6cYYykfBwyfzimVFCjHL4e2
wiy2Tjm3DSwW51zt16GgZN+KIx5dv8eB6R4DrZel7ogjDpZ6exchSVww7Ob7A51ukKHGmLE1py6z
FGytmITwrbUNjY3MWgNG3WBHSwod7mtA9a2mpLn6WppsJ2eyw20XtQTDj+13HOGmPqh8qpiLRMGv
YuEeBZklHtFpI0PeE5BiysrqiedbpJeXeZh3seBLo/msrJE9vZEiIyQxu0di26ucgThlTSRDo1HF
Q9Y+jh5hg8lXhWsB3Jp/Rv8tVJ38iiVcUo59n2fCpFW+Zsq24jn8q+Qda0W0pGafUytBxl97wCzH
/vmE4GOzwcDMJyXsRVLa0cAVAiCLJMywOT3JTRppWToNmWLBSBXz0Thrjsa3QuiURicMLc8S7sJH
eTKECVm8yHm6ZNN5rHGcX14AcOSb4tsksRuJh2x4zfQ8vazuQWfTTjs/IbVr2NT0wYhYFo8VsaL4
Zuoc1zkTsOW4D9omHCUAMTfWnHq7MFJ7a1W/ZMElNkZ4A2nzLkR2S2YCwjKd0HB8ub/+eVSa/nPd
P3xzjhUfFKb9L/Fn5f6OSBhbPnTo4/CE5sROLKBy3yfNda/u5yFxkyfgs1YWMelPX1V2Ed35DLY8
yH/Xn1Eb1xfiPYqt80V5tBIiOEvX3h3Nd3rD3wKaPnfqfhzqQAuWRO9NXMn/FTqCBEpYuSMG8ybB
+21CnuWj+Fx96FQhYk8yF/tD3m4GEZuT0aGVQ3luiQeUndt34DuE6iTAK5on1u2TFt+FT+tgH9YR
+xq8hhJcU6o9ftOn12NBtekSobNFoWYF4zjfXxzzxlQ6ca/1KFl4q2HQLgAnItXSvXapYQls72F0
o+RF9xl8DHUel1iXwKrG2DYOcFENLbigdNPkj7EObVVPaW26N/qRT51U091LgWc6LjEJM9Uz+J/P
Su3l2vVXLX/PIuTUrjzyNJ2f1gU/vrhAkygNm+rwZb298e5oukoBH6E+g9OUvDcTdXOTk4J0+rkq
KmzcVdYHFP9TjLtvOXmWWvcVVh8th60Ck8XzjZLWevDHxGZx83yHwSiZK6HwextcP91hNtxJMiHj
6VFQ/aiCnCI45PA+q615nJO5mh+NoJZrrZNAjK2IcSJMUGDek7NQ7ZXgORljSnB14WxPQeDbAfuN
hS9Th8oXxk2DyhDXPSGLrPRZnVfTLgDtXjalOew43Fne5V2s22Gv0CsHoJJPRkZQrmuJPfuWdQXl
P+Do3zjg4J5qgkpdnPEusZzfAWruSokEFxvn3sSRDk9ffW7pxRxN677pPkVY1cXcDH+YMrt+Th0X
Figuxtu0kCvUt3G6EnueNlWi3f+06Ul5X+OlR/VaExgkAB8Am7KkQF1azz9hHrf4mp6VtplcSoiB
+GUvpp8i648Qi2qEQ+cx9M4QfRrldDC/FWNVm5wq+OKLF7KTTpeH2d9HFUm/QEi26qgNOHqbJzy0
0PW/ZO5bIoIzcnEMFwLYBrRJmmMgTKzKds7fXBiNfS39MHHeVs3uyXO9+7TyjQtirBvOQloTevxS
CYzR1gVPF13wC1uUQv7olEwJfsmKR4x/5ODttWugjyQz19adtUaeEklETO5tnAORg6957BCgoE5M
n6G8Hyaf/41yvoeTID9VmLCIH9vgj4SUgB36Y+q9RHWEr7bJhf8vQVAgL0gcJOnfOZ2689V+5vTS
1gmHawMAZGI57414hYKr1E4ymGFe8+KQeVYxQZyI8ARDXG4T2WlH58Ag78+ETTdGyQttZBlNASs8
LRvLAE4wYK+WmI2Hh87KBaU9YT67BEZJ7ErTEg3OqRUZvVnaHYx6baJIiEZqi8I8ZfzB0F4GsAQp
qOUcdft0g4OoD35glAC1K0q913gMQ1XDkgzXXO4HOfbTDsXEq9DrjoOBFVlNIZX46NHRfUDXh8bw
62R9KQ8Fh61l8V3VHGoxDVPTJcOLcxAKrFCep76I1c1Sze0Q3GOnYiPYI1ZIWcDyUhFjZ5R6qR4a
CFFKq0mtxIY6UAloSS9MBdYsX21VGr4FLmB3ozpzimL8CWQUhF6/aGqsXrGOqn0D5pz7HRZ3MKG1
ZRlBHSImAYwF4mnVcwVLCfrYrAVVCbfxhollFfBPzyXW4cS3gzVSJrIHvHt2Eu1cUa8THpdArchH
5Jr5qtspUwmfsq9X3co8OFj9cFJcKnN7YaYKOhepbJQr+JRNHosY09B+L5mr6V4zCr2bDpXmOmwS
g7xdpU0Utb55OaFZ4keDyM0cj3kl29AMR3ZeDTQHi5zMbOJ9hrPeDIrjVBhsl2gEYhNfnUsD4JQV
C9EWxsN1U8IS86QEFns3sxQrcWPk5mRfCj21IQP5anthAi55xTdkUBQoThHntnRWFxRseHBOvvO5
p6p2PyqzXzZq39ivEcpPOHzr7r7gajzHUDKiqFb3MOV8Om8akY9qordAx+EQ1OWZtUU4Q9twneYB
PhhR6GiNUTeK3TFFLMIjoRATFYBgOB4IK8tgSCaXHLD+Wit2Bf+Z1JRsS/e9MlxcyPCZV+YR6iCZ
k/Kkn3ghl7aZ7ncST9b43PHMkYvexf4Q7RQKUnX0O3xj/KCd3XkJwxb8M6flZYSgwNiZLfkImRnw
98lq1c0lrhFNOOcfcEKn+3aHZRIcPQkO878pq8ca0NaosxaVKo/Qbpjz7v/Sa0TD/l5BPjXnQHDV
jcW6wjBvB9v3WjAYjeV/4S3aQPdnEv3wo+LNXIecfQbOEyaZsKXU4konJTp5RCKSghyCUZJ8keK2
VeQGYJf0Y9zRcX23H94YpNZ5DtaATb+R1nEpMjj7+AeVmkf02fQkNzxnebHYhBV4DKRymFaqAc+k
6amueOK7qhs9pN2X0UcLblEnJf7WwQ7W5qhuJlyyfuEP7zhSXiaDtyOXGSXnro0EZe3TuX5I4/m1
JJoGn/uA83a6vVNyfdMbENVNsttjZZqluIfS5tP2xJy3grq7SiBIdW7pg+ic7jA0LDwEG3Uc7kSe
E0GPH5LZlw0ZTZZgaVv3efSrg8sVDyvk6pIoKOZTRy3BnFqVneJUxqi0WYDB3EWcXlRetE+sZqMb
AR8vALC390IZdYuc0veoXinTUCACnuV6aI+8CBUVzlUillHZ7P9g6FqwbF3+r/oIA3RathhmF55X
z6/Joy3RHrL/NHG4oqiN/j0a6lDdvkMKcU85Ied7Q03p+YjzEjj7qdCZYY/iSk1miEhORS8StFjx
DBDiVhGWNig/IIGBNN4QHVA7Qk98kM3jtpr+iAASZuADB65bh7MYuWroCvjN5NEa2lub8yRxSakW
VKnWOXMdlvAUMrGRq8468wVkRbdmGmtdkZGojrZYh9LzbqW1FjU5cJLDul2iRBSvMPJXZlsafMZi
k2B2pmUXnB2TtYwiaAd0VACWDa5PRo5CRjZ34bHHIkpMQuv9HwZAzZoghhdBNXaHZj4cAlRFYfFu
Fmo8+FADV3MJapfzZ7BAq61+m4sy0NjauFzJXWBk7YXkRAw7KUvtXIKNds4KTQm+Cm7CrRu3BIHV
97lQQ5eXvLJwAJ+VTFdQLSuCJozec4ERsq4pff6PYNhAYpULj0t9MApSMDQWnH4bw//ZYyWz0ZgS
fDhXd1ubueXH7G/18iQzmbwBc8qZayvFEFI1iIbcdiTs5Q+nSyJ911GxlwCF/S7B3xQh1Jwxlwre
rP4NK5vYj9tw07VLI4LHCbwDZg3hyk+kQJ53hEuzjGhO8Gz/Tl2X8WHbiXUkztBv/NMpz8pmzRbi
Zyk5o6r8U+Mv2aUxys+Ch4sR+gA6u8BjgOk7QPfh4s5p7bTLC+Do2a3AMIkV/4PZ60pnAJ5Lkafl
vVlMQHfU4aOmIBRoHKyp/4EuCrjrf6XeO07gKbo9Q/EP0HT3K8nTF39cu5jOdweAGJtJmBVZ1rNL
DOWffBH4WtBcaGkunCjcQsAR3uE3yQB228iQltWyIbaUhCsPOmOP0UgwlhIQuqO+uKS/553t4nJf
2SK7/mDP1RLAVt7MM7peu1qkMYVsiqCJGMhOBGtjIsHCcnQS8d+iZcrV1XAaff12Lika6gAP48fO
9WF8HEJKrve09fp1g2wDlMcUCZqaFRhRs1IpRf6pKKnwMCkoIkdg+In/+O1s6LozVfsqR1Ngke05
fAP7HVOdMfsW4PNLyedTZvPYyLRJOOMDnkLpuKxHuQOKWbODp95A9WavAUdz5hZNYEgtgTkQ714l
L2O+WbIxKllq34u6yYnJraYGvl+VM6Gxi0VHpSbWTha9czdN1Uteuj6fdSiLXJva2Zx42Ux6Lpil
JbyGV62wPwJUFbearQhx2E1H47G1L73VuEv8yFpYE2FCcpe+PO9m+BbkFvELBmxsRIC4GD5b2dnw
k2JqqDgXac4HoBNSztnTJhODUYLKyuiQFwH+vjz+q4V1pca1S3Euf2HWRVQDLarg6D9xD3QQKqDM
vm3RaLrldgCY+1F5g4n/ucbYvsRCsBxP+XQmxap3wF2z8bQDCvNO/g4BsqAiL4oVsF/N4/5OzRvI
Ef4sVlWvYy1EJWszX4MM4LC9k0hhWB5YdHlduOc1ExGe4pS+cUdw4hLW8V9QqhitT7ne3obZKTRd
Xfk9e01ud3QmeSW8RULxqxiRb2xH3Z6nYnvf2iC3YYHHSvh0krP49ybhCQDeGHN/yvo61nLQXGpe
iN7gUYiKT0oripUNOC2RKqwzwGf1sPrjXX4eR/VCg0f9xX1Nom3FftTXQWhlqwwXBlQoXNMNtLqv
LOxMB3duStJhAfB9GFofUTK6fWy3Fk81B7ly8g+tSxiNSGFNUu5RSj6BLJUoYmL/aH2ZrzoPWIWf
mJzn2tuLjqK1gdRoBy0I561nECn51zafNyv6fHI0ntcsUPsGHybhIxeQ5shsRkmPgxsqKNpcvQuU
eQeVV/Rv3P1u3pKEvtaFWw7DIEzbOkau60NFuDuNNYcFN7/W371TNI+DGag5SvgMSflYT+blDyA2
s00m6nnxABD0iiM0msYVqDqQGi50gb2Ys3igqrqjhi5zWKoQ80oXpFU0cnaI0/N7ujk1atJ7YvPK
ew/O2+UJtb1Rxvr55To6WhnITontf8I2MUvLBaDOCWbFQP3tlSgfT1/d0rmDE+nrPzwC1DxNjHOh
fXrxC1faFiChekdJqQKZqp9rsAUeVo7/mOr9nO4UinXrvLllco/mDKqudZy6wH986iFuTszJbwrN
m34nd5/XyqjkMft47h6hyp9dyheJhUOiEIeFJkRIYOG/gA4ApYmBZOaOY/XO58cWgU2amGtrQBvH
iddnk/XqgCI1LA0H7nTr1VtZCYLPDZpA0kEJx4lcxQHiAjxaiUYAIKmcHcWHHwe7yeN1MKSYertY
fSG7FTU72YsBVFxyMD0CXtW+HC0jzCpbWNiWs1sQk7JiuoQLi5w63loCy9mdSU14t/WsRWnJDyf9
CO9MDtMF7tcXv+z368aBakFUEFfQ3qknFZSFLYwunKQvnII/+ME/CCQ8epOaTDyZVwARy4dPPfMo
szapLU+lTshrYRspdGa3G8aB+mDVKZwTKSz9IroqJmbA8n8w7W4ixoMrXOiRn3nSch3Pbd4polTE
4ig3dPiHFzPkZbOM+RywhGIqp7ORVZVNV4YaeFpWimw0Nxyy0ylHndlVIxES39tZ3x83brkiRKRg
VkM/ZfJuL2oyIX/D89JQHcwt+w+tl5tipONSmjMG1In10Qi8igGsV59xUEezoLg/j9RA40JzyKrV
4vtXk53Z6Hp0p/+nrxs/zuLzJBEYDYqQx1AUUgaTuTCbFqNqav+TuXlzFKxx4kUCOU3BGFzK2+1z
B1HgoBZyz66LJQyjfChZCmgUtSDTOXoBuhzcgZb+iIzMpc7QOZCntWL+RcbXmQIhIQss/jFz4daq
sBKBj1kbh7u52dUsNvyLiUhTmurQ4gn8R3x6AVv6iOGJS8QsCdav0loMLxwOjMhKgjXiLFnv/XYx
Bp4v5pepqzvICaOYHqcozpzVSmKZ13aYyRbMSOVClg+5Y9BLxQfTCFtxvbbHBIQEWo9eIyPrIueu
UC0m8YqbjXd3MsuOSM0QSXwTFFVT3bCFWdd6p5S1fxiD6n239mnvpFgLcQYbcXBayUTzTU/dTQrI
St7UfKU/7a4s0TXVQtX/pm3rs28z4jnEED8tN6ybFr/wc3BaXUNLcsaHg/KH5SsYykdCbMLalRkT
M8UmWjbL09nNzGLVHr5SNHW4wudMpA19vIU4Q0RiDQI8UaFXw5wCR+zFjQ/6qLhN30SGXEntkTME
WE0FQZao/dLuGtjZBy1ibxRMCbwwRy1axYhHIPepnJ6GaqeolhMfNJd8E9j2Va9oGEPdriALhjdI
3xUlN31ulu4YgubzD3RMF4fQICtq34r9HEkjT+MbJBeu/sRdFRl+4Z9+yHWPRiaGfJGVPy50zvCG
5HaktQ4zu8HenHmWnMM9h2C/U/RVZ148lCoaX78qpy5x6oO4cgY5n0j/3pC6h8rpwxdRkmTUftJN
mBI/n2FmpVvNNKpvu4zllzBygXkQwEp1hdfxRtp/VJ0fQwGilMlQLQ7ShfXRq04Bw0l5ItijWWst
sK+m2rpeOUGpp0xCDkjnp0+dvLZIZTLe91veJHQyOGjt8j7fO7tOqv5XcDMRjj5CGILHp6Qb0rmm
jAsS1eJZ9rwQV/heQONqJqviNKQ+xYkUGN1C6YnrDDtzyf/hUmQw7o3dW93/1xTB9Vp2Sjl+OcGe
5z7dZs2AGpFh4eP3Jy3JJHQN05SodP+lRqGMAntvMqejARJmwJ3mWMAnkewBVEPFDUvw5pPoOCby
Zg8++jhcGvBWhwOh74wD8l1J/sPG78cxE3jh97jKMC958FwNCEEF2m1aAjc0Ma1z4PFJPwWuHv8V
j2dIdYi87osUmugeh29t6Z6+E4G62ZgRvouKqBTKYFPUf/jGtvWzw592XIuBEcf+i0V8naEWierN
ef3ChSq/v8Tq9yQ1ONdMYxa+WSvcL7usxX/FtuZSUdcUrVZJG+Cs+D/xksCTvGW0BdkcSRL7O/8P
eCNq6Pu1Y2oOEUIDV5L5oIAZEQn0VQepgMzxqm5/fxqOFJ9VtKnR0MPe4dsed08cH6xoUZVyQIlx
SuyH5Okp0RqljMMgF9AXxmZp07FApmkDYksi1p7L1vMW0dRK4d2Z1zs5ZXB1kvP85tJnwy3VXxro
2wvXQIR42JDqVZxdZV8gWjtAIDuKntZQCK054ltCYMoQzuHPJDB4yP5mI/O+owcZm2Iyi0I+704B
Ufh3BFUok1QDROlc8Zzi2GpJYBhMsOY/kTGp5h/4+2tVqk5PBdvxKsxbSohOc5xy1tBtv2xMtOU6
rsbfiA5SAZFb9pIcKU0e1n7qGL19ovlnWlKNzmeTeNdughxSyAD40FD9iiyVs8Nq9GXBtwJvzGq6
for7OEqvDD4+DI97zNvy+lMZxRCEKmJs7GtqYCsiBCQu57dg843/lfVpa8ZgirVxtROEn/XGItVW
w4dps1U4M86FTMoe0ok4ymrwjzqI4OMD/uBfqvZ1zOw58zbmzCPDVvs6mdGxak/ap1kyBUwmPCA0
PHgioJtWORnClWe1h+JKFGpapXdMrKNui4Nqif00TQ5gUh6Alg7/0xrqN0TOaB8Xplze/ysfeC9f
0DINX4Ph2PNxWn4Em9TA0zgyxuIbwq3H2JU0rw+lCV7N/L1YLgc0IdHMVYU5xxyqIiuSqi0GiOfZ
A3BmVnrzXIPkJ+XP4YdUJzc7GLACXE1uRV0O9yVR8ApDOs+grV0Yfp8e/+SyvO/9LqZUz7HtT/GE
TyuyTo3XW9Bh7SYGk6ApXI08QIUUqXKqmXxAf2y7lHWjrGxX1ysw0Grr+KEEnbayKPGsTDvkDu+r
zdE/0uAdVhTighFCwsbNzBR1Q+9xXBdjQr3T+HKcQp2ITHj75/u3zJg2I7M3cGmJNcPX8gaSCvfd
y8xQqtHdisihq0C42P1RlAuPK1yLcsq7R1O4/2FKyhd/4cN0FJlPKBgAn9hRA0gWRryPrRjHykji
j3nErtYpMzG5d099HRwBakgaEt6cKKZazW49wEwIU9vfxSz4zNgXpg+1wnUZHchnjM7VzLltG+zw
AJP+LY7kqledWPDAg5sNGFdUcmfzX4fx0Fn1GGlfvvZXVsLxwtboo5GZ+P0lXg5cGVkxvmevjpBB
fPVzg0Fq07aJKXiHllAIEtZkZBJK0xhQ4B5AfbQ3a0X3wbBjrditFGWdhtVChwHSM9w8YRhh8jE/
XPdoMEIMsD3vATGk3mjVdQtTUO7JDcM3bxLDWo9EUzzPEXbBemjgvUY4VaYlRmQRH/6fieqwe7Yn
TlDxz//kh/ZJXGbJnLoFJLl0mh/G3RY789qJAdQpfgQGLHl8k1ii3MvvmcyuwRGhJrpG8S2Pl+gI
Jpqo55JggpLgORpc6dmr/YPKPPxUav1q6dkwOz3xr4L6yTw8L3FKEL72ClT9201TmeyBEfD4eISO
L0pDNJ9jdCxC75jLOKulD0phM51qR+/9Wp0pBuJhKHr1m5ngo3jrV0Hhb6ZWEmODwibrYQH0oFF8
eN/+3oFyqJr99DFZcDHOsmHbUeQ3eZeROJmTTKuY1c3o32Vfoz/1NFZG8LpqeifFjHj5frxjb6Qr
2Fb9eTnfJYcV2LKKNCKDAgOPKOUXbAs68mEHKGj0r0L8GM9it9AfvPsiWn5bLHSStidoxt1sb414
KDr7trZ8l+EGQ8qLk8SsHm05AY80avfDu8DHrj7alzh2mKNp7xftDPd9J5b9RcVu/i9484UR411r
KD4EWPjDeNR16MZw+7VGvefSfncCoystxSwUk1bbHVReqoIkcgMtozh+ZXQiixHQAaJTkfHW3g2w
Wk4t5IGATQwwpe3Btlbqn62VufWI6wNei2pt8NVpTK8GKWQZK4nviYLPjax4tNSiqV/Toxda+8d2
TRH25FG5zIrlOCXmOZcKuHGanVeN/YstF8pSgAO3TC/JK3Tl/ehF9aEO6/iy60G5Riwnoae0vXVx
5VMe4EmO1FsuZu5NyOYPYJuqr6a5xMhUo5HfQmDPKXsL23szxSvC2Q7fEQ22+37BF3s0SlGZ8ysi
K36qZ1jjdF35/hacqey/vsg2PQ+YHm7w6MWuTHelcL1NEv+mAqTvjPAy4W2gqf+5i6YjxltuVDXs
PBnFNH4G8qdN0ujQ44U7qk+NXEa26c8eXx4yj1OM7qMQwQjotvCJamC7X+mpJEjI4IdOlJ7MAMVc
6hjVsyAsrK4gBj+hY/kwnajIutdC53Hb2GSwr9Hrw4CvhwQthzNQY1AhQsDE+Q7/NxeUUwpuTR6o
C7mpMQiv6a5rZ/2BEw4YuV+lJHZCo4kYH8onVabHiehg4517RvuRt9L626QUHqAaxq6Eh5a7Bzv9
fymHzooFbSjKsiRkBi5SAujI+Lo23w5T5DwpRgeN4qlEUreUZVJ8oqVO6Q2C+sa8ZuPvrSi1ytwc
Rwh9nnCQWafE9PCee9U52MU9/EHJVfMARYwj9IVDvSL2GtLKWRbv8kmmzcVgj+0MOWxwVKPzI9ys
oMVTeBPnjwHHIuJj0DWC9HK6Jem2MKDzL2byVfzcH25WweT9AmgSCu9hVJhstw/gBPpnPjccb65f
3PvIYEuCLyAYL4G5fSqlFqkHzO4lR8kMwTuLXr0Pj//231oBO+lDeGVkX7V75cGKkmItwh+xhLTR
hdpPo93/O1jkw1CDbvLHzIoCI3u26ZBzSozXl3brIcUx+yYxvw6zTTN+mBbr9IkC/A5bpt1grlF9
xsK7XuWiAireEzDBy5KewlXhsS8mW13m5tNMWhja0x9sGv5IE4+m5TQ1ZVSp2KJRi5jelTfP39bt
DbzAQBsesj9ERMb/k5qmanthfskQhyBLnI7WWl8Qp81zv3+r3wivsNwi1Ny4/mhoqMjLbNF4iAdU
Mdh3etTVkcM48ovqi4uAB0LtmlN+cA2u2Aan6krVn0YQ8hWPV0l1DqrQj7uiCxzqUEtAj6No7LlE
MY56njlWOtU5yt07X56RAagDMLxNntGFlz9xyoTAH0YPskz810kl2IkV0DXz+9dtC7Wo0ZqdOjgz
MMpUckmWJf/xmkxGqGKbJ6zotc8CkYO38uBjCxzfkOEBNjxNrTUnby4H1ZGR6nryfn+EtA3ACtMb
BO1/1//LtZ5Uun5u1jyW7eRm8qGdvvJ9QqC+cIRGvRhktdcjLW7c2+NkWbUlOaRZuMIqjxbbg0ic
VDuqNyU1KHs8EiH/AXvpLHa3yT8JKXlLUUGk0NfpfL+wT9WHPb+g3ItjUz1/K6DEHyDo5bFcTHDb
xMsuZkDLRpGxpCinBZha6iN4OnEFSuvBEyF/4Acm2Uk1Tu+T/vySUvozGXOmkuuLBwou9i69znaV
aDwbYEhJOUViTCnOIWM3XtJnukQg4suEz0NXlR888L0R1hdBSsFVJ0YRWxX70UmjfVFtGCFYthQn
yHYc7l2/3T1kKiQmA695knp/zYrSw2yOkM+9sLCzm+l9k0NnGz1w366jKce2zIO0zVUjsSPSgtcU
nqq3JiJJIhHL+muaIm2FISoqoGlk2TQTZT3w4lFceSOUu6RK2FjY7qJJBfRFSj78qjInst8J9PwG
3Hlde/vN6j0SUgwt8wtBpuJRi1v/UrB5so7/0JF3R77feU+QeKz/LCgi4PiEMD/i0wKFMAMesXa6
l7BOXmte+lUnl8xAIuTWey3picaSg1iF+pi9NgquXTzUVnyrX01GV3NB1oXBiA9qB5En30Zkut7g
lXDYaNOkxf4ZiYMc8C1k9TC/4FhAa4vJn8gqHODUegTGVzBU+smPsdLwOZSedT+UaDlMFidN21ZK
3BG/t6Q+0s72fp9ZRQxvNw4AHikz0UZH8uqzFbQ3y0Bb1WzRXPwZ7WtN9FjRXreKI46YHGkRNdLc
VHD7NMtZxNqmFyZ/x4OZrs3VXMdquZIceZacPH2CeFYUhKh9TkxonQNDr4AOjzgrBfFqoY1ab8a4
Po4Fx/b5GoBC5g/gZVvk4Zkoaa5nzFGcwoVn1H7gyfwHnUTxNxsyFZnAcuKtiL1dXEQL5Um8Q6Jg
OtEC1QlGlQChvRoDiHhx9IDxtyrhDYvW01ZW/ub47xlEgLAmlACbX7YQlvy4bOsp2Mx2t/66+lu4
KFSZPE9dDjgB4UZJqK6OFGrvd7FXsPCzaHNFi5REAeo8VmIwccmGP31N6V/FAjRqdGAzVV7UVMsf
RIU5DLNFi3iLWr3YOI773ZHxjRjM8YT190NCX8in3/lvSbDWNN0FJzMTy5k6SSWNRp5Wb4qG7ez/
++uJvDbxcMWxg+zjeX3Zj0jj5eqOhd+Rq7zj4+h1N64kH9RC9RSSQi3ju3S0015hHZL6v14Wp2RG
hWldSLn5h63J4sDTP71obe1ILyM3UMow8GMlhXJgbff6wnvVNRZwKeGg3vLDwrahNN6mcyy9jlT+
v1VQz0W5seYmJ3hPYfgl66Gp2y0gh1gpM2ImgeMijgvwGiyVnuJtiTZ5U2Hm6l3v3urU4hvqp3az
LqY736IfiACGfNepz/l85qQJKZ/OogCmjkvd1HN9tV3oHv6ZugeL0unJPEyBv3UWi+EMOX1+rdA0
KMiXQRHznzbSf6HuoEPXVlRxbNkMlYJ+lroWaBJjYdOdZ29En9nXGqyxIpdaNn2WHhNRf3dMHFwW
6PP9GvZy1UV+HeYVq6RGLO18tLo+LSok5HBq4oR6hvMCUr4r2Xn2EPaIz4ICcYKTCkd+TPujN9/M
iF1lBE8Xie5n8+TrEy4tup3qRjV7ro6QifYNmBxPkj0F/HQB1v+SK409+c//pp/pArLmqQLLPevR
o/5Q61rS9GaUxeaMRlw1PLADmYUw14WmBjyp2avCryk5Ci6eTIkj4AZrWpo+0Dibfn2rR/TNrURX
zMtjRePRg722+o4n7A1Ja1H7+ZdBNfW2EcCFql3QvehANJ1WHedU352mmb/6/7IixMiNoPoj81Mn
Ow6aZtABo6+xNbZKxO80EKZ/rEEJ/dMtY1V5F04iD8VDZdQ5T6dqk3v5xMpojRNISpz4TlpmeOel
ZehiGt9rQgAuJ+eoG4zBtZCNpPScNQzWQWTE4a3wU8dK4UmwllYWa+j7KsJeWb/f1VTJ839LVPaW
Z34lqqwcfvUZnyCNXX3Xugfptrn9rp+uki+JjwjJe6X5aU6mROgt+Ye+nL9G5SG/1OFXZbsPkKpT
ABxchhwgMhnnvexvWsMwoX8Ezryt5nU5faN+jKqO7Xp61aX+uRl++csrzQeeSvllFLIaf252K6g/
6s4WGWszYIjeMNY4QPvmziLeF9f5J7An2cGEeFQOuTDw5Rk7c8vaoL5PtcocqLVywsgOIi70cqLj
qtoKS0mBP7817AeL0/rDi3bzJQvZmtUbw9xU9G+bQTzI5sOEnRvPT6MaH9cvxo/vWrHaiLgl9Q3f
EZgdPtukgy2W4YSmV5wYkn3DTZfgNP0BXu8UEMj7R0kiMlkhPlKP4hdcO1KhoyZq/fkVXJ76u5tu
ZLpBtMr1CpQyydL132ToOeATzuhaZ+kAZPotiKtFgmHmPVTa1VJ5LF/OC0L6izqHmAhJzseJpg8v
pX9K89qQO0EXbolFnZrR/C0BfXzsBpaO/2fMtIWTPuUO6i/GufYFSN/zmioNvlLjxzWUhW0xnHSk
4cAltaTUFtNKL0D7mSK9oRmbVR0lZXlxWnsd5FSOCOC9a9Pi3BvR8/KzwSYSStJy4Nz8IG0xXEXH
Mb2lou+o9ycB6ZYUMAwWTTF77ZW7Add95kEz3sztV7HJTX5joy+kw+a3PQWFBGRMRX9CDJ7JH71x
Oc9F2jHpaNllgSkh6E1IR4IWEF4Jb/LIALUkjwY7fUO9hpMBn3jqAIja/SDDOg4naJRb02FlR2uN
kk7Uqt/I42r00r2Det3f742NVDSDTrm4Z9zm06P+5dN5aotzDPmYD1ubqh3ou4de+05Uj0OjApLF
2NzVIytfqlSacqD1/UA5xS3RuI3bkpqq7TD+qhYhZGekbUNObJw8baJkdKnNK1YdNJBon0F/A9Xs
G2ZJWHf7+RoXDrBjbMIXb0DwH/917D/7C9Ckr7GiZxGwkGM+NdO1cTdT2qQhEiqjbmVZfjjN7AM2
vn+PyvRNdp4uurMSuKNKRNDVf4/nC3mS6Cuw2nGFEMcPNET71FQ4WC/c4rVhXuhx7yn6C4KpxT7Y
Q/dwP5T/Y+8CB4ZS4hVwsJ94Of0VKLvCOPDTkdfpyfxKslbxGoYcZis/wZAKQ8xXyi4E9oY7swtm
H9Wlu2i8B8+1Ija/2Se58LEELVjGm2yedl1vx82yURwWBbeMvEhUNytXWAzgEZR0BEr2H5ALlw3s
fKhIpvXGakDvkGZg+D9+YWMVKQv7NK/uUt/NVeunvFubAuuMPVUFKE4wTALVnDz4+iPC51X+R24S
x7zrTU3YlxkdW3CQ2QhcC+s2he3gRPxdV0h65XfxuRhJwB87Z14zc83C8LcZ2hN4rBn9Rs+0tTaH
WmNVWF1eiHGoK7Yde2aGfAz8RTZS8meh2kBtI2a6TFLbNajjW5kVh8PN2i2x7wKbGURjN2gtW4qD
wa0t1jfgAkaZAEZrmfJsOqwzFmCGQjbmegxITtm1RmhaZPUgmFQCRlDdSHo/5fP0I8ZPeIEAG662
KlGlmAdj2GhFA9y2tInu+UbrRuDWmqQHLBz1eOBNdDu5EREMg2wwI4E8kFiDbKdDqicTldyP+6g5
gyjVH213Oij9XMEJ3B1ZZ7rkEhIA6B1FDDAKsNwFd/VC1253XBxAN4Eu1bREtscIZ13lAKilFYGs
l3b2YdNNY0CUV3jOhBUSG8Jf1xKGKCMFwpNQ5zI2ejnleWngMP8JX8v+Q9Ij2hLLiwulyedRW+am
gwwVu9cwyUjW1QWM94kWcHDQlpC8zhz4/JqgGQcllkSbxXr0ksB+q6VW9oNMGOKRbHn8dtqFD4Tf
u0hBGdAe+aKmUdiOnNrXal4rmJQsoX0tnNm65IWcJ07Wnqr41bxSnLUnoP6lkp0qWU07ATh3Qf9n
cLWLojgzASGIr2fmkqUiQWBpecG6i9ce1WtBENUs3R0iNiVvxhBHswRbtO6mPLit0ccI0EKPh7JM
US/XNjKSO3akghs9vjzNJetdsvSVV0nuKTy4xiITPzejbPO5FZ1jmLIe0GgFoJ5oqdgqtL906d07
tnPxmosT2R9BtZ3otkMPtzrl1OYpWTFbKWarnilhfVfeIx5x1rXMU4jM4Q+wDLU2qkoVrBbyxCiX
MZ3aXrKHo3NQ43sXE6e+PzDidZoDn2Twq0lprzJCqn22LazqxDnOiS3jgh3pIstVPIQkmGFzZ3JM
I9hCccrLdVyy/9Vys2u9VXy5ZpNvCaPbQDfBemEc5CKhdt3hE8B1B1cRmKv2d3mtbtOHUxehvRUi
Zi/7jr3A3ahGmVe/TvRRVFk78En6JxN3gDKT2ZCuWgptZkspHSj6VspbUUs7TAFd+AsMcM4BSfvI
n+xyk4Rm2065oB/KjGeRJlnxD73MRBTeRBsL9p3tTZSeBgtcHJhfwLoJPpDKfe8TLYmOcGLKp5K1
oi2GgDCetsFLxy07mdw1GrhoRS0txuVJFswPcGfuSkWSFHdfhvbpK6K+Z0DRT1rjwvTyHqSMXqUA
l+lntHrxCSr5EJL4skk4bzSsfseilKocwz79pvaJ0/Z1abqq89EPhyNLY4mBbxsCo+462NMG/jv6
XeoYPFCoDC6MrP4CAcv6VzXCSc8a+ssfvM1H/ACvil8Iu29wwD0Iioa97PNkSRAL3jBCQwlUrA7m
0ujFxhr8rMvjai351r/fjY2zYOcmhUc8nOSEpGuFgU+Lzqzi2KlvgDzzjlHLr73M9f+F5yL/4cbS
2wUAX3EoLQhw20zpLHz9qXNEy24XUbr+BWft9Wp9JYgjiMyL58wl/xSBHmLXO0MPyOprRlGh98gS
0HK1T/cSNZ4M/92+cmobGUPTNUbbD/PRivBcmvDkeOccUhdowHyaGoFniBPgnI8z/fyZ8jztTztu
fBzrNutkiywRG5LdGL8lMqM9rOZZOxoJ0PbfLXt0G2kbxVuedX/5qazRreTyZQyXfvpN8DBT52Gs
i0l6VDSKVZZlL8P2iqKSw3lz/+fNKjxQIlnVuZdBTGLdNhliMXrSVbAOu7bEV13lxyjgVrQqgFiW
6xvw8l4Hx9WnsckRTdRvRdgnQ43G/9s5UhQalD+WI2uEi/sZeLxQ5no2RLH65fiHZ5j3pQCyaNFG
rkcg0G0hacx5tWvK3iRaY1SrAb18ZpHM8+wFsp2ghcXPIg2JYvND9u6dPWuOWyIq3TlheVq2z7+R
vFWZu+bj7aQ2TqjH91srzrpEJzsIlck9IbJb8sxnMUz9Ng5kM3dJifwQwPnWlQvm5GAGrNV+2BB7
AWW89xgTfst9tFr9JIVztHb78NvGICFhnQrhOQCBbmzqHmC8myeGc/B26BfmY4A4D2W0k3M3GlSl
za/bum9i8BJ4Sqz6JNrU6a4UwPqLXGUipB8F9WRbxCN0DJSepagnLiVjRH9rNiwC4R9Y50huCgxp
Sc9MjONAjkt3g2A92uVZuTWeavRMES26/F0ytnoUp/7nlcowctXLmy5iHfTPojz4eVMUyqWYcT6e
i77dALZZ2vg8NFW/aa/dPiKnve4iwKdcfOQ3iGZRnRlZukmkrRPlnk9GxTEItViGbbB/HRc1Fjje
/ndf6+Vf45rY5Jkqk87Za+Y5CRKKkxYWBybzRIOtI2EcU+fSZLQRkcl258wSaijowS12BR+rTZpj
V7dYodBSVrmg8bUFgtTOz9aaZmpCCTFBd2hTajyRDRmOMl9w8n4LyA7uOfPpY4scS19xRFTKlDq8
P4TCI7HCWolVfwzAEM52yKW6EMc1XSXqU2+NWOeocqZQUq38F4EiqtNiIqzRkoPbePQbsrF7Lc39
m4FCa2MBof0TJFnoARxCbxH67PF6vDqwGpXhf005qxfHnabBXJOSKcAgQAFOJLaBT6reJ3wUPnI1
mbneERYUW6oXeor8pmUoXNUf9daiaAc9vswUTu+iXb2Z31iZ1DeIVy+gSMI+a0LSzs9Qo4oZJuYf
39lRaoXHOWeWOkSPJLEKBcw6D2ffGenZPao9xJOuYgXhA+y0kkvIqYkSKIQSYWdMA4XSuUyhv4Fc
TtPyp3EoqshHj5UxFwm57Vy8xmlHQ8mOH7XNbWqvmICj7i7PoBfW13NvugoiE8GXKiZaMYueGQLH
QbQ8ONAhb/p1vCV9LFjg50Hc3lqiFLjrjaCFbQ79xJ8T59kZZFTmYgSy21mmcACdUMZQFFAzFYSg
ReuIOj/6V1sujNkrNxSvuWt5gUfeoHAr6ogQ3TzOVMmfJ58KEeQWGfw5MZLNwWyadPDZ+tkVWlXS
PcuTujy34hmt1tCiGfGS7Qv//8dl84OiaDo/19VOEFFCYXDRvaDqB86RtX98CE2ESzZtXWKFGGb8
Fi+j9kvUBWqZVULR9i4VZI48kneqN89cdlucIjmABPPIrXwefgRjPYo0MvfBLh6ffqxanEfQza8D
FUxPayXNyAS+fcFqPnnJEGEL1DAwJRyHtlt8BmeJ+GW8XTDwdWoVMfjyUywLabx3TgPLSiD+AEF/
jezN8nG7Nl7eblimsMi+DdOEZIrNNOUWQ2/TaAQC9VTEuLLVPCwrENfnTlqzFGn55D5F8w27J15T
kMd2PMelZ6cgrFSL93lDkf5+RLsaqjf5JfTPt4iaKkaHivthR7ohIM/R8uY85Xx7Oc3h2MFeoSNp
otWSsbMgaJutzT+s4VGlXaYXT3ijccr64FzAWKiogdpQsJd/olQ/5IoHZ7v1XgbeJFHGSEhAQbFj
7sbz1e0MSu7eUkUx5bMPDOj29QMp20xIsTdgQfqRMefkvzGS5b3abkA0mvsNqH8uKVOdGtapLp04
1GUexYU+ovdJbocGh0yrnKXptFVvYeDsWbV1/uR9YXGeBTHr2YbpOgipiDFFODHxfaNXZ7dtKNEQ
TV5upIeH3IydqWDvdIBTxtpaZWLkezuInxeSjBpYcOJAZqlOdqyfn9KYMnWuB8aepi0aLw41O42y
mSUhSR2NlnaHtuIZQLEC/sIJ5JZrxwNX6fB33kMKXySCTH3B/aDS9dAhwLx+sfkondw6HS57qTPV
bCHT8x88Hh34pklyjZ8DC5uxhbcmxPRTJ5SH3O72Dk0i26dBU4fpbF37TXQIvZywIDeVqBqXIWYr
0Gt4HMa1ZO3O5aWcIAk35B4HBYixGw0T4HYRVgrboeqYm0kLi9/783/ZGkW/cjqLtUZjEgv/I1ix
Y3kwgQUvxCrzqbWYQI856FTXid0VR+DigbEoihT2K4XqcDN/fxjZWbV7ws4ajqs6vpniCnIfPMWV
eN6lUoGzjnyI7GyvQ7qXmuDbmFUtoSLB9OP9rsjUjO4sL9g3wtJySHsxLkfjXiLM55A3q+Wk42FD
wu2WYhsvN8YWLwRYIaIyRryKwEmLRucAI/YysUVHhY71Ae7fCWS/x4gwKJhGOuVc+4eimcBOdUNS
XjsN1gwITqWsTsarUMyJr27Lq/xGZRABUwBD4nZ2hPENVf9xJjCMmOEyjwC6Give9EoUpGgCJQ3X
2XUniprktUy3JUx4e04I77htmjnwrJVwMtNNRrJ8t3y7mYY1lDplv3J//hg9gB66bUdeNc7XBf++
S2Yl9i8v77bmx3G6qaEY/UMkJ6qNq4+ehjq09EbirBGayPIm1bTo3BI5bWAcRia5/4eAYgnYJkBR
hWGUnycCvTNaL7Arh5rSP1P04r2WT33OObI19dYeQBSNdMwmp0YRMEdkT2NTR+mJHYaRFjBAuaP9
sr7GHdyGxQFGrwciIHrT4r/d06/pUrSJbBp2Js25qEflUxFyuj4v02RcoFRXlF/6+Ny60X1Q0Cvb
m5V0uVWfZo+3rZHLeBkFqqxrb2o/UmAYhdspsToGWCMXibxrjwnLyVj0Ybh77IRvZOTCK1w/3Jlj
p8owrewEP4B6P1xMXd1EIV8vocYQ11NFoJMYkgnZ1ExMnFOt5NYTqVpACJQt/n/ipPlyA+r1gaX5
/g6QHHblolQbrSDbMpJa0Vb07EG64Xu+1hYf5JTMvwsE5OfCenVjh7OIH9r0+QYSQe9i6JazHIkV
AWVqsOqwSU8gMeaFudgXm3d75mtnzL0OJfb9hFfw581tFv6PQhrgiXPj7vGIAGUwf9i5ZrkYDzoD
3jQdOyO1IH5obj8hZD6CtMMczA9sdCAN4t5kQse5nbRZvYRebjGK2QVBT58Ch0ClYjMXogATdFbH
WCvpBzt7j4EwpWBci9UmrJp3cCrRFAzmMgPt0Zz/8MYjegm3uKd+K2hOKGTID6vmtWW6gOZJ1DCW
jTQDjq3ClbZdQ9kyN8N3KQ9HOx696L/dFscWgJw2vAow9jo57HVPo+XAGP9+bNr+IpNh9rwGeDwW
8o1MOzORsLgBW+8yXkbBT4+F4cIDSwZaLht/aZiVmFRhqsZQWF3QBGKihU5cYeOZJIQI2NngSZwB
36ttVf3t97ncLA27NYG5O7F4xleoBkFEfNiddhGqYjBVSBleYexEabFNVbXTMP3zReN6jm0yDNEJ
c+yBHZeKr/4qq2WxKBVM2wOdz6JlctRLKuqyxT0GhISZ+KRPW+zcdZnChXC0w9PoA7x95AGemImG
DUb9rMUE1g29MhuOQTXvtfmdsZXOuN0PRYlc9nDHtNyVlD4nHFm+uxelHrD1hByey3+rDCbHZfmx
ie0h2jyDIoS785PTS0wsyR+RJDTNiSY58fv2HzP5c+mtHPqxxBFCQHlHnSApiYBSUYGR8ekVQENv
T43Oc4P5ijLFx9IyDY3NdwzdzmBMCwPnWNiYy/f3cldmw7NF5zvj173f+T2PALYzhZdQRkoVGZU9
Fy70+ZmVL0EZafNMPT8tqIBVvi1juFPDm/HjJblAXYj9ew4ue10me5X0kQd7UKZsfvTfR25DFZpk
dhg2t7n3/gn+LCvar9y8dUIQ93JDb2jRUkQLYurODAj86K+omM4OBhiHBQupqvnuNcSFw29bYgvV
iRdayZoAwSkqGxhkhwXrrMQftvWAe8aTmJnMLt+WlJ4ADPxNXOW52GOLAmhsRIF+1sthQ1dINb7C
yckWaMcvRqXocMMDQ1a/2AhV1BkOAHDSK+G+PwlUp1CX01c7HXvs1d1ZIoOueS3zncOHS/yUiYx7
41Abv8yMJektG0Upi4mtfOCgffYGp9fT4qsGmtJEayBr1h4+Ib4RmiUh/KCwqJFwvfCPBPq3lQki
Rm2zKwsLDYRqk1kwjTegvsCGzB/2VjxVNbPAG/OBkugT+D4f0zXs3hT+G7qDky76y0nCR4oSPNxR
M/58P+0D971nP9Xofrn346B7EVeJMRZq8efcNntJdLZ3ZwlYfGQ6nfO19VfzoC78ujkcgvT22HeB
HW6LJfHdryC3gWUjBUcJ/6ANmrBjvGsiWS1/UISc7N9DpKmMV60bFeBMyDV8ontMwZX8X3u4OChY
N/xby5dM3sjhBBGvHmrzRpvsS2T9rxIR3HqDcmgDej/Dp4l5moAGAAG7LJ6RWhYQPbmefccgLqAI
+sCIqfVWSNn6uDWJK4uHO4uHIThFoR2saHMmXeARpttiS1nJNA2CT/xsCb7g0NwWlz3bIEX/Ki2E
2nNKXhXJUUuFRPcTaVVue/xY/8dENCodd8PHADXIxzarofTZgu/MYhQnK8747/xWhvdJTNDKknKo
4Lgzjmk9aUT0CA/xg4HqNjFYMVoMLtp6aRihkXVNMb7Tjpe4qXsqTUFd7IYNIS+sscjJf7YZPh00
Uvrc1U/o7spl4N+zrpkAr4xm09yUSvkqj0n5eT4xVU3laKEH4Ku61/kmJYJnQi5HbBKj415HtTZd
jveqAegSSuP95tUwAprJIJ3P2rMDWPcUMeng44NVj3oBmR6gTyM0DF/VWaHmc2FVIL7cdagKpMrO
Nbw9hXBzx2RLZjd82kPFWjbRQEozaHCaoxCWeO0k8ZaXDWV4/8j48AValUBuISp5d9HA9iv608fl
xk5nEwyA1zUn0nvRyKiyksBvepKfCHJTRL/e99DIsJzr3fVczjmVX31PPVwdfKdyFlQquu2dTuPZ
TX6og43EWGKntCTKbsq7aYl1CkgwwQLNrmaY81stHNTWmL5q6KMZSVNL+cQrQ3jERRozFOhCKhLY
1vGBftA8IGiJTyykp/sRFJCrqAltLG3i03xr/2223AUSYABbhqH4RVxFZw9LIFvVUp5rdyAHj6cz
wjt92QzsXiuBEvdhnETmcgg3NpRKFb6SEhwT2ib6Nga1qeMP6dmGz0J+GqLZz91u/nj+tUoaNnr7
n9Hr6gcQZ0KFFkhVhckY9vs9gZ5ylTwe52QtIuni7LJLtQXrCnOP+D/8kHgxjTuXQAA1+riZNdh2
jNTnCiK3uTC15jwE/O4ThYwRXrjk05/CjKyGaWX4r9au4wRrGiDsHM3X1wATDiFS7HFAh64SzsWL
vYq5kP5SYiM1Zj0XUOOV34B2TS1rJv7fTT/NfzBSaGgKYoKXGsQSlGV8nnMMdD0BDeP/4hB3M9fm
zibHqAgr+ClHhCjqmO+k5KCn3JViBYOWwnL8hutTzbX47Nv2+IFuuSD8DAJz3T35hUynx7JajSY2
sRoUIUYGTmAsqNII9UIqclxwPELMsxWWx6RYpKQem7i1/fFNgvOJGGlFG5fHuG/Cgx9AuSs1hepj
vkSU7jFb196Ma3XYdHZB5Sz49qs7Mr3LDaNp5z9ZxhxQXyOD9gFEyc5HpQEy0NkmLNK+h7Nunkv1
YyAhC0NwZqcph7re4M//I4scwl2GK2//nM0hi7mfaj2EQya2c7qS6Q7j/6sD9pRhR7O+m50vlD1B
Q0icZDV1n0SXvl1MWqnF3CXBs0HPUF/QjeLGedlUUAFaNV40IwXsPx11enioETRBocWyv+HaHZel
OorH6xOcTESOF7al8GSvuRPuva4Sg9NlakCdk/31fWyLT6w2HZpchvR4sGjCbJXl7CSRgNAQa2jS
UhamCWevgzljbGvEPAwCmL4aUDSG+i7r4KKL5Dji2C7Rn6ZNiHsukf13rHyXzxgPbCc/TkdlUp5c
YIFULhtvfW4cVHSfdLozoAawekOH71R0027JqfTndcfK+ed4YjzpwgpbU1EHAjlabvYSaBW8Zq3u
ZjyDMRx/LGZKmichAgE3ZelvInDKDug+IY3K2HZEN4ttaXyOO1uV+x6VNNyyN87NB7/vzcgXTb48
JbHE506hcr94ud/sLuv+Y35i/W0IvVJ4d2zoyz0pj17DgWVzxWhNPmYNYtU5s7uEDJ3SBYpp1WOb
VV67JQTJizvOiUJhbTVDmkmXsxY3Jkq90qGPsf3ntD3Y//W+Lzz983Uymv/U3ICqSXGpTdRsVg/H
Negrpgu/xIRkyCZ2XUtD5KxbCcaAARGZZV04HbWulKJbKGASAsJczgH9PY+N5EOhIBSwpD9RfeVq
pKniW/d/EJfJTC6jWZbh1l2xZKVmjweEaa1ew793jniG5SxMdps2ypbK6ea5SEvI7UPeAIn3Ya1x
APeezQHNpA036s0tBOvtMSAqGTjKRd0gsIJF//r+/FRfDVY7wUOC9Gw5boAoQK/p9fBq3NpfMECI
0pia0mUvuNFI26coVi7BVrosRLanqeGpN6ull+NEvV8OsZri/6nWQqECA07q4184gfJmt8nvlLtM
ZFOlGw/NWDWB+9et+SdV/BRckkh48sJ0JdmRmAw4nLyytV1R78z+9u6qQQ2IPC51W/W/D1XTIMox
jyRTz/IHIokLRVbnyTaXKfKfeXhojYZd3PO5LEUCrw5eJHGV4nqTi0QT2cWuKVuqY01V/Mly6ZRh
AcdsFmRe/VXKsmmTS34KyzRIWr90KCTlseszCTdcHCkf1tfUvQQDF9GZ4efLDEwOLQIuuAmS5bwu
Li9JQjChW34+Yjyg+LN1gldjmasSRI0E+hm7a59Id4/Vv1T2HSedFvC9yDAnryHwePqjwFuOK3SN
mWk+KU6gIKtmtd9E4AQJTmAVlW0xsvm3/9pNoXynA3N3Eagy4E+KUKAUdCUkBUXlH/pQFSgqvy8g
/9/beLmjmeTk8zXWKTxyV7BTq2PB6xjUKNjC8erzdbUSshnh/3jIW3oXNva4y0W5zifyEc0ShGWV
4/tD204oO7iZ8jEXHcsJ82PH6hUy5mFn1ov1Y9uo1/zTSKE4/y0aZZeDm10oIo1pdqQZGpvsOS4S
cp6P8SR78JHOAPqIrQnrwEheSMfRebPxRl/TXRDY0Sv18TLS8ZcypZ+qAAPPNb7OFkvg6VwXbJzQ
Fl/IUH7Od+DnlhB5mnSp3jauCH8fTzIEWLzWuotmp25L5BTWXCHPUd1TIXhFCb/C2CsRyOZGdNCm
N6T5CUyaBLpGTcuCj3dPw5QicmnONqUkeBS7NJV/7w69vGA43ZQArTLpDGJluuHFc9r8fnRsJzCr
Kvhre1QkKcZ3LY+gbvsgrmMexOki9NW09kOFNXOSiCNapanCW2p6dzSF2Rco8kcTTx9k0laFFGeI
6o0b4JoAAYcUmEJUHO9+YKSJ7L4RXJkth3RP8OXbHtBgHbCJy5y774RQPTXhSGk7HMJF5uTieaqA
kocP+AzR1IE7HhouhEOK+F2CClz4ZOu2vHdkWJhV/8iFB9S0aFX2hLrIq+20WEZFXGv+qOheMTsm
JcQL8TILeyXzw55CHErEhxQKqpj2mEEJU53B3e4Ghyk7nyGixANllDyJsZOkPuVO/vCOMyhb9NT2
mfJ85dJuqRjWT5e/HBiJoPPlHXiELlWDzCv0DhYS7eo1bsCq9H14mruAa88J0bKlr60Agk87uTJZ
5bg4fSz2aLWYin8izB1oCj3zf6IJ0l8W1DGS1sVAjzS8UAWmZM6O0EPQxi8RscjXlQwIP4GRdp23
kK7+a4JfLVqMH/4Sf4W7ct+z9Wlv8p4c4AOMKzKo/96uyIBYYk75xqQERL1ExyrYrmPuNDcB7yfr
+B2YqorHy5VdxtNgiJJ1BwuybsNRZ8RIy/OHkPyfyTuRC5yiFmXQZEOyjGTuZD0wG6SMalCWb4rh
B2p5EZHF8netBue4zzx1d19riaYYA/ib5S0ZHXR5G7E+mWTK0SinjQVXUTdxZC+c6zm42odSWnkj
f4Pbc3dr43igC4H6PnKLQ2jqeGRMFDfFhf6qr8vjDT2IkvJR2lcf2BxM6ijRR2jmQUpYq2RtLBGc
++8KrP95p5qCc6DgsrMu9LPAYXOjI6sUXtNcZ5F4xfJK9WTBOro+9egM1IAv65LS7Q+fSKp9oCZi
l/vde5acnY0sNW9ZenpAl+6+LzVPYT3c8Ft/ovfznMe6SFRDAnnzT8YpJOEF00P8MBw92NBWhrhl
ElV1UD5HW5BXiLBS04JaCXHpqjggjvwjX9FGfrAM3MbMmp9Sab7mY17r2Jvn4tv79ryszNz0f/hK
rL+ovahnqhkaHxhNEikPIByUWBn5/W6+Gi9r8WkEXIB2WroQVRfLxFZuLCF3Y3ZwRvaUe3B+10f9
LwKGzcFU0LDJJd040tZSpFfZs3/PraJ4Qj5SQZ/Hgc3e6YgNiNiPhY3rdzG7bYU5scevL3KwSB0/
GIXjDg2AogXCnM3n+YE0nCgn0jeFIPOOMu3FxZzQ3fMv1GmwkRSY/LoTWDXhJK9If7kRoZudJHWi
dHW4XFzPvb0lqelkB4xRWA61wqHazOeu/MfTedDImFdhJDB3DV7xNFACgci9ULo7CWd6E0WhZR9+
3gj7AKPEJ+zPnCm/OGQUPTwqjLX8kuaIqJLqyBiMKoWFtP2ELOhnwvZ0cMuL+GIjtzEbEnsJ+NSZ
an4xjDM9YaIunP7tB0UTr5qVBNkGVb5zFDFPOegft0GGr6Zxda+14G4pzCUeag9zajJMgwZtxHox
1XbUMOajDn7twQdqpxDYe60+it/rBuXVXEBRbevAnk42YRxDfgbIdEvUZ69foqVdrXGVbkIS8Mk+
CvuvgAJFYuASZKbhU/CNdJlt7OXFhYqb5aDURIrd6Umykdm8H+9ZY2iTcHnjBNHGw71dIZKZcZx9
OwGyRfDjJ85n701Y52e3tPBrZyGmjLvAwjmDRXpNEqSDout2gI3Mv/1R2i7rEVnfBjyt2WPjdFm1
lVLaFJk3iCyGkmXqbyZfFsZCklbx516KUg/epWypy3ZW8pAN0CX7DRvpDcP8uUU8K1tRLa6F1lHA
8JaF1UdQJQ+xYNUGIjDvrtTSE9Q4EApX1qKYvCnjuoI0EsQRMXcNzDOGcW0VDw7oDSdj7OUboBc5
ouOM4jmqyyer+Y9nGJoOQF3ZPcpa+Y8ct/kfoe4udQs941B3Zu095NwXHPWoWSwgKS16xvUAPv+N
uPB3rH8qMI6N2K5dr0mkp4ZYOXmjNvOfXqi334E6KD2IX23sjERFQ9zisL5+2ZdAwD89eDLSENmd
LZ6R6e0GsFLCXcgad5hTB72xkZtEeMUpvtShgRylOuOiJxgKL4cSURKs9AJQv/Exk5DjgqETN4/T
YojNh7kDYI39mfjP6fklaQvrDgg6VedRpgGn1nc0Tm1i27uLtVuBDFY6OvNAacpdBh5FqYm6vIr/
RphAHhuq6QAQuH+IULNn74t2oLJB8Vz92Pg3if+iElLLjGDfEoAbArKP90SIt9ULliowBUqzkBus
4MVcnaCbRiIEft4gdmqFx5cDwSfObcLZkcbmAp8xA1MnWo3uhs3qwDCWwdscud2gEhwCjMF6euSn
KGMHI5hQOZJo2moNYkIPQbJ/ifMaYC443BAm7re72NsZ65qDGFjWt0nwGbd5uJsgnu1BnlgPj42d
dmqISLAtjFE1KUtP01rCpPOewSIlXDVFJmsoTm6ibKcKd0AnKC1IZPAo3Di4/r5iQKk5Ka5v0Gsf
EgE91RCG+4+csIdGrqV0ORmMCPFjVTjieeeXr6cCOEdta3Z4g3d4U2rJV3V84aNkc9tbdUgVJe8Q
dkYi4h3GZ+TAPllDhz5+dq2eElXfS2NaFZ3M37bcSQV2oArbTLVBW+dxz61mIP3GHLf40qgD/4MN
/Pa2eBoDsA5JR0Oimk2X/JUieV0bGWHKEZ0yFiLcu2dwzrVu9MOFUse0I/k5ExTwqD9ChMau1UTW
C+hyJ+puJRqez7KGlOSgthDMg9g30MPMUvqtTnijgGQkCBOJAqxzhv3U1Okqssa7MC4mRBSH9/B8
bEI9x2ErnH8Y6YygxEl5IlQLeVk+40o1GhojlSEYJmTTNi7ym7NV1NXkNsRY8fZT8D/xx8MUVlhb
7AymPj8fbH0qlIxVhq2887k4OFKrmmZzDlAxyBV0hLcOP8IwlrSk7b5fbBPrWwO91+1Dq2d/1pae
nWUwLX74AhBKf0Ktl3z2XVG7FnL4DG3oru2xPVAPrIsgo9Gpt15dFdSJLEKYRqANCbw/sluh79vw
yUCvQyreYoTN/SrOII2Iz8FEq6tGcLb/ps1w4R3OvOHI0dWNUg75es+RAVML/3+P/yBzW35kip5M
GVxYp4SRqCzTbOYuC5q0t6wyuI0a7vGEFlHZNXRRB4CpI9teQGUnXV0u5+kLkiQGNAIWUVxyHO/A
uUqRDdXMWt0AI6MvYUrcZ1ILBysrOaWsBtal+IfvJeHSG/ms/HPT3UoGV49fWI4lcKWxHTWh16a/
heZhbiS9HOfgDQ2/jHOaXBCbKtp9vBJpdBC4LFynLsw3d8bzzKw8QjWofvgOqr+b2QKPxaBIiYQH
BKBPlPkN9rryCUQbJa8L3szAKsMH8ew9V2BjGpCgru3k/OS2lazRKPmzDWnyfoZMe79TzPQ4t6c2
GH6V1fpjz9U9ypfZjazbpdIAAK3Omg8eLiefqBR0qsTKFcOQEZlRPJyORTaD6MWILBITVUz0JGqp
8hd3r/IwEaYje8MMd6zIfLHi8f3mWbR7YQO8xml3enrwX+ElPs3SRsR67m5dPKdRx7qUGGp2xsfK
ijaM6jlAdWxQNHjd9HJkPo+OGWJVt0kGKlRB+FUToHXfO7FGSeMIX5riMksSXfH5yx5bFS20IaLW
p6XejpMdruWsRJjw2yumz5ChPZHoWdw5ItcyPqnKdg3gWjcJ7+Ndwi8IFsgN7YMBgKpgF3xhUME0
MrMVWCBUkORLu9dJQWdsQ3/54BaSLmoqikgSdiv2LlEECCdU5H7lCN7a6ab7Z2aU9/M1zQXUSD8k
ecWsqrfTZWtUOIVnc8QGYjcvWP1KCN9cMCMrVCCpogcke7W4KMU5cNwUMrI7vMkSGDDUgOzoLASQ
X283pRbhPQWbMjwm93AHjgoNcZyD+7h/BxI7pcL6wScMm0XYEMWbBQw9+kyNFdzCl3y8XylQaYpa
R7QECWlLTczs+mD9ZlcdG3nE+Zl+jfod2RAgWeQwhIz/In73UPZiO+rMl0Z11MJ9fDPETjBUy4bC
/DAPaanxQHrI/KjWhaLVQr0uNEtsOrYruYAoFY8q9gKJaAmULQIGeau/uDOdfIo7jwu8/0H6wami
OkOQtTrqf5IO7Tiz3aO/CYwpXNJYSf4PAbpBZDkx+CBJbzDmTaVkFbURU/yHpIy3RHVo4S5NeHde
Xeyr8Hg+32EgW4ReY7iR5LJLzB1n4BGvRXavMHzaZn04rFBf78wzYVthBr5LJk572cXF6504f+tz
hSAk5M0CxYV6e1hVfPvc/msGiW56wVuwTOTpsgjOgR7Rvuk/EBo0opVJD/KeIcdVB6qn25GbqrJC
18Zqxn/XVkBXcY17qOnZU0ZAMZG9DLhSl9/baAaW09WW6f4GRDyIL+cE0Xl9XHP50kEXRQ3mCRPe
91nmxEhlN9aBcF9SLXcxmFfEKo8F8htvkSapF99HDcFP3XIx+ssyVwMLuDjCXDuU+O6HvsQiuSoG
68/MCf3PPzAUKIWTqtV/XhGAAn8OeZFi9wTaP55pgg9Ki3WJ0GoJHGBZi8kWnR/hPD9fKQWsx5OH
ZHs74f6e9cTJMEjJZuN1z97rF/NgPXKGmJb2zWMbErTmcyiQaZ2CdRJ9ukeFJRrBRgIpJYoYhlsK
kfHDA/xYGuliGQUI/Bay4wdV8muzR7vr/KNezOlXII8hmr0u8XrD9uhHpgnTAWBhdfXR8KWuzJEu
Qt7lZfFuIfxVOZ2eYTVOPrvQlFezFUBQUgPb+RbzKyWM5G8d5LCyNytWGyvU54MGOgg+zHbz1FI7
DQugIo54Aa2SjZQH6j47LVwg6lGssnq6Y1ieu7Z3KHhyTIjPAYjE6/FjfFHrGwgk4PZX0/0TgJZG
KWE4lIJL/I5xLKjmwBYkeMy+0e36WgpPkKncPlIFhPSzppxEHP+d2UPcgr33Wppf0MvaoRTLtN0C
1abyXhDYU9Txt94s1dbHfvsfl/yUvvA6Xx9SDwbBDLUiw4cAkA5iQwQlKIq/BBnDZm4o41RWriMg
HqSzkzrGkTXbHCor/luV1NKWZ993terK8z0l151hwaLGASWWsTnKzz0i25FO3NkHaUoktWQT8W8P
LPk0Ktq9uqj7ZMuJnuUyyljjVfHmh4RDcFnfcUAigyKsQHb7D7PF5Bl8lP3Arln5rfzLQpwghPo0
m6/lA1R5zff81Pzt+5iRuZzqmGp8NNC/G8cfNrwNBUVpQKxzT3NCChlYjJ3Wv5v04wrhOySb6Rdh
Ik6j1g5/hf5AQ1fvuBMJGedhaxcupkfkkoXuecDOt1FkraAuDB4tGtX75baHboEuBaJ//+o6Q5Cy
L9VI1MTPiBeEg5E88JeM+EkyRUpygu5T6RSmpqI5BwRa9PryyKJO4GWKoBdRZQmP98C6wpQkkZZR
nMv0mObRelvedlqbyp9TP70F/e3AjP9vpkiNWCab1yxiCNPGynEnlll6pkSd5l7xfHWbAiVDpfd+
L/rR66duVJC6WFh8aHgnqYE4An+TsDqXzvTQmS1K7Rl29nzEoCix5HMkVcAO2Km8PToBvGrP4qPY
YBDKfuS7+wIHxngtNm2Tsva3OOAAd0RqCT3Ler0S1JD8DVSleZ2jnTutWRvWX4Lvq5i4v+J9FlOI
r2b+2NuK5A0hlN6R4J8+///MUArTnSciUkLe7f1Sdn2MyUwUs/K9dGnbhtI1vsP2JrlrQNPgFsIH
sK2218EzBu0a1mzWdJ8n5n1ytoKPFNi7GrZdQtxYvrw/MFafJlLM99CPqroE9fqAbaZEdg6EaA0s
+PSul2l9qdsgu5XcuhZudJansViAL2AMczQbvNnpJ6T4lPxzAFiLvmwYZo2WqVueNTOtmdwGApq/
OjB+6XQfTN3vQJ+X411kMaKuZAxsQ5MoFXsinrkyns9N+z9rRhW8mzaoJ6vpGh4z3MVY9BM+k7hu
yo2T8pOXtMbdHBf4ameAsEYQFmCrk24eJq2Z+RIx81PfQyHq3k/ok6FjPKk5B/kAsTfYmBpT2/3b
8FrROAenDIFbPBB0R8EGpfD+h5iqj1wa/3ZK8mGNY1rF/L5EXWjet5YRLeKHdVYQ3o0yomo16t5D
Dpbz2653Xn7MpuP04i+HBjf+1xvCyTXoptYDrf8CMqD7+FoeZ9+PJy3Yyj15DC1+NAlSqJDYhaDo
emlFFjg6TbAKp67NhYG0LE85DAGYgWAURzI8spxn6ZI77gbC5gUVMUc9YLkYZpxQlp5VP/mGDdFV
GQ+Dcc+Atho1QRDCz6WIKNij3MKD37PyBRW5jv3R/vz6kGF2/ym0BzQYTRrRbZjKH7DnJjpOSFTO
fMRE5oTZztyt5UFrgy9QIdLCvXLsSyOrq5D7UYVF0MRBVEdkbNP/ivfQclvuNsCSfwqxvyX26tuy
1jAyc9FQTlPm2h8yb/SSb0UAL0tBJwuLT8UXNdeZDi8D238BewLFVuMAfC0uYpVcgHIPGD5zKyQ4
WoYYVo5dH9NfxM2Djx4scwDfRP9o+DEQnw293A3GrhhcjyGD3+bUt2+dvyR26hG1JcPtMseYqYUz
IjDBvzT53f5jV8XRCqbr0ikJl295bKsFy7ddT8HWB/yF1dpxwwOXTZd5qt0rZFT34xqRgsy8kVHd
nxIsTCxli2HiI7lsnEnA+iVjIwTA+6orUaezuaaeiz6tkFvzDZlSdLXo0P6m9AZfdr8BLqZxRZUy
rkvep6d27XkfkFrwCHcMZ6jsdLqdqfLx4yjELm3Z4G+kylyF4ioK8ZHNNATORcRPyJ/y85aikRtP
y0GpN0TG1EAMANmS6znf/skxmnGDhl+YkeHFb7fuH9Mh4noq3ws1REtHngplzTNXwC/1exC3onTj
Ob/LjSJSwpePHu3ZyIH9vPbZIGSL4wnjs8rvHiIgmwmbt6LrjUugVnm6UmjBBLT5S0xykd8qkyQA
A2U5l781pp6E6nTqTPKUP6FFak07GwQl52pehS5+ggStFePHTOKiEFgR+KH+uNtTxnkTrTM+Ib+o
JHE3i0BY5MRhZ5j+sHfHkeW3HlNkYKbP8XaKFQqNrmhrRhjPqO9e6+Sj3ePZ3JqnXNamZ7ThqYh3
qEKktoWhyGVH8uZ4LlIPD1OEX+3E77V1pYZEim+geJR3QibDjgfmGlM13CcfUo33fP3nPNGaIjNk
62c+76pcLAflhIB3XpRvv2hNn6rgq5ubKTbjx7ZCVmtkuWYVGFMLuYjrh9FX08pcLQkPrd9+fhQO
MGM+fYTLBUi0naPTuiTysbjynb+5rojlQ9LQfVPztaniLuBXSbm0BsvAmQDOEf+pKsMO/mkXXowL
e66barftw2FRGvBTWteQzRp6s4Juc570S/WLve1SiYNYpSKlRF9juHR4XeNg6/mmaaYU1Qx2J/9b
qfq4aaJOY93tBfFMjGpId6i9kDI1FtVwixVE3nog8wlbGWNHOJa+pNMLBP+bA4XRE6USvAGaoqpF
KyRCda515w8jvWz/RMZHPlL16oFV/tnKpg9pLLV9jJQH62eTuCBmpD7He23NzWJiVXXN0Jek1HT5
EDnjEjc89obEDlqWe+hcPoDhjgCc9vaR2blDW48kclfXiC/SYPG72xujn3JkOIbcWLKxfNUvjMmr
x8TXTGsL92dCTq5G0sweJmWNHgu+9GImGjCHf6jTj2gcsFX8jtIU+jV2sE6oWFghmyMwF0Lo8KxC
6fAazWSEXnqdOL4o9/5PVNwZiUSDu/7Z38M+n8I7fcdJebTjQEhS+RrIoiDiD5daVsaVOqY9MYSY
Ney3+/v29l5NubX5BzWw8mulKLYHOL/K0c84LmVcU1y4Q+m3G//FM0RNTjgQaAOzQ41swSRgsFCB
g0RvQzryBrbCUWl3ZoSoHb2XasoNn81saSnFE1yO+UmnWRO1gUZtwHvztjAyVlBFG7pJm6a8As8s
3bCzznXf/nisGrBps4hACGffelqjQRY17mHlPl06mJ/3QDsuPdJzWHBG2J/Di8lBJ/dw16CGE24d
NHJblBCL/15aIQUP+Ccb6HSMskxz9My7tp31NLR2DaVA1sP6oprejlskYlMJUEq2T6BMPnVrr/uz
6UNyMmqWFMhcLG+iyS+RMlOzjKeiGkA3qNsiRX+z8V9MUEZgR2Rc1ksuzmYb5GW11jZAMRTdpw8X
Lmv68dIbQXNecHoFCF5bCnYztl0lwyKF4JBNVmjsg6/V0fMqQgGXKcrhJqRXimMZVObdCxK+eqZe
3Hj7KKYU7Un7KWkAYDMfxE8B5aLShMzmg/OcRjMmCyBe3QmocO9CrecdNOl4nsXVuuiQDeGMgn+1
fF0DJGDaRBzUPc1LCEmuc9u2JRWCWu7EImOcFtf47kMNBit90LmoH4Le4aOmJ2vgETESQgVWSLb7
6G0nx7SlHNkb2nBQ+x6vCq+qrAcAWDxm/U21OSIufa70xoSUeZMFMenPfmHcV68GLY54VLpf4B2A
sJAmNUJCjJQbYannrlcUC2WbVDlbM+TzxR2RuOwCpJzlgltEj7O7tfc2TGVm6LOsaB5KVl1HL1RH
gpNi3h8pcCAC4gkErfx805eQOJFsQxWYHmAp5oJ5xUhwo30m1LoqS76mVzCEDNd4Od2jDt1Uylve
2RAk1D4vzwmrdAlK7yrjXIbRNraMFHs993CeUxCFAc1NyJf6cC8S0BLqy4fHEd7pOyH5c/gNKDTG
SYzJTsZtN1EDptZMNpoJNFV+G8k7JRh37mTBdu/SvXIqNoXmqggfxu2l8WpPOFQ9dEPSTWzKFyhS
uEQxvM2JV9HFLhMJEGU24X8IfFJseGXZywhpcftWX9FQSOYpS3eyMu6DhjxVZBYxvGGll2zfkIoU
U8ei6MGmPoFlgB9cJK7/IrZCEcZBQuvshy07qYWQ6jsFD4WfIlMB7mvTHrYeimlMOMrlhnWOVSIK
rSEt0yj1AnANMsadLz5vWS6fCy088kAzkscU74Rw6gAP5eHWh1OVUpCWvE5Zlx/a5ijGshrJt7Nc
KbFfx7w5MA2CIMYP9x8hF5p5oLe2fNIIQjMkbcSuRPk5MTPGaaO008abkw376Q+ZkDSIBj+ayPRj
VfjBCZb/T3ou9vmWhBlFZwIDwewdh//KC4Ujw5JlMVfyJs9NHGxyG8dNP69Mxrr3MqVUs3Ooq8AJ
cC4bqDYEmuuPrdXCemuD9j5fx6WjWmQaoIZg9jxttmTyjUTZFFVvJx3JEkVYyYcfSlE/6jeI3zo7
MW1UJvjv9YZigYU3Q/BB4X6rMFA4JRaJiLGzs37TV4CLa6Q6Lrnc/qABflndBirFcr+JXZPjitdr
BOzKJp7Dnv4+7LBamvh4psR99tWoUKhIKtGeWN96yHYIFRx8hQgL5Uqt3sSeQ2oGRCeFyIdCQ9Uz
sm5Y3Kl7t8rTtw9y7ugDZEn3XROt5vcpuiW9gQDTaIsMommro49vVU23OjxZIB5cgUUxZWgMcj3i
grtpB/j4N1PoNiP6Bk1Z2FuyHQgd6Zsn8i1aCYgSfO53ISX+JgwNsiGkDdAKewMLZth53MugPZyN
sheeJaEDRqhq5A8cYpJvm6rqIJ/Sw40sOr8OZr8EeYPQdEKXz/PV/dJBsR87FZGiLlOOqCSyZqgl
wtkrQ/SOBVXAoJ24mnHC/dnmIC5O6lkiNHbfhtZraSd4Vnf6HhYy0ezB5gAVMrZVK2djjt4POLvl
0TkG/dS5bAqGXkQBoUeFpTV/PdLOxDEdTiiNRez0aJhUfvHHgc4sY4nodK8CryO/7c01uKsg5ZHc
/s/7IU15YK09rE8z1pS/7YzLUGLC2+QFxHaCmFOWAmfsWiJ8gdORcQYCEcEi85ZB1fCgLEDHIaRB
d4mgd7Ho0OByRFRyh4WWUYoNdfLKt8XzO8263beiogvFxSfWdkqGEdlAVO3of4E7MsEUD8BG/2lu
RdFEiPAqrfux6MmkeHrhVPYArVrrWRV/ILkY2iOpZJ/UVDSfB0SyYAXlZI6GE0N12amh1ZnHUxQD
QLf/LwGD1/BkFwAOYqwrfQntukSQ6hcBRbECw4Oc7fs+9RPtxynVncDB0G1ws6RCF9Zmn24/2gXD
t24awiIfUutZr23KVQiRE/BaHsa839+8GoXHnK/6AV5JgDpAcTQObIvqEwHH3J9546F4DRCPX7Cp
xBGHiteD6vPg/KpJIYIhaoKBIkfoXfJsDJmtkK7zCdOZwM4NOim5ZLlK0RDxB1uEx0qQxEoOxLjT
Cd96Meq+QutSmm61eBHm8HM4phlW+fZxgeGj7/3ROm/qgd2BLJTDWGVRk2juokO/vqR1b/QTTSKt
O6ySkjW9aL0FP+pVOmfyHLLTYL7+nT6aupqF+scg2yUl7kQFxEScSc8oKlziqfCtwqzJhWRqy/uZ
wlM1LNY+FyV80oDYLJ4W+V0+TzPycyUPb0jVJURTSZK2DA6HejLEXIpRrhrp62eDeoYIk9TwbdcG
vI/fT3MeHbaw9KFav9zTmHGV1tE1myYjOYITotcfZXF+oC5oJNHG+EiBjI8DNK9SqFy3T2QDxKsZ
CsJAHZBl57Lh3JJ1Jij/aL8/uDU6RV5D8lL6sIdE5fjHeWUkcRuIV622ON5FprEJzzHWPn5TZWm3
Uhy4Ty59+ljxV1lRP4a2l8Mom95R07tFldHgX3deqQndpqE3TNN2aUKwu/LJ8CzoyMLmQOkxwCrb
dNFLQEEjcjss2HM3EtHLa7NL5EHRn6fP/jcks+d1Pym/RRFDr05dzGxzvlna22bjMUMRcdi0otEI
sEVPot7OG58OjvmL79pBOcnC6KcK1do24NmaeFfDiK1wRV3TDVHYX5S7zp84XMc2pQZea1fck609
u2/1XwuXBXNaH5B5vvQ+Hi3un3yH8vp4MRkXn8G6nOgONvbFXi7m96MPWrs0LZWUtpdgR7hwz8N4
fp1p1DTMwsIrKRejkFSyVVNiPgmqKBMlNiWrkKjgaApZHlxE0uwXzJI3HKprbPUFeX7XwuG8j2VW
bcMoYfVxsVhYvhMObf0kAnnK0I6oWR40c0jv3AFP+jtl80R/TkQWCHHTpjpFu7D6JRRWzo0swxvG
Mztt+T07AMLogh+VCN1iHObReFkQFS3/DbqMk25Z1G8We5IFTu+BLhhkuceqfzsDmD3tjmdxq1li
6NAtdZ9ru34A9rCTULmrwdrSAmL0hu/IK58F5YfGNVM96/5kbgwvFUEYaL/UlVV4n5YHL5zIndQH
DPsyyVXg001xbF1wcNQlDD8FUM/pGdP4H7dEsh+CRHPp3joOj4ms4CKy4NTioMuVJ7TDwL54DsMf
hiKwZm1ZMNEg2GtFRqLiDqfpX3FqHebqXY6qAEi/UmMf8jhV2gjoYI+MklQgSwYdVivasuhvHzfe
mBmJNJNG82i2xdmAdXwFiFRHUdsd4wuXstYwy7Z64Nt8Tc2zBbtzVAKoLaGACa3aHefzt69IMc/8
wLgOsE2W0V5Stq/2FH2/ftlSOoLBwqbCPmj8wSb3YipYtQOplhC2Nb43TO+7R8Nl8NSqHD7kSBwF
/E5BYcESnlZ7+iVTu5vrRBlYkB+NoqfiTdFZv7fLh7ftT/B9WzJlFCJZQ+FSmhnLwJExLtcOHa0l
Ap4B7u1Jdro6M3EOc9oFPbX0vosAsTLYc95ELSuzE2meaYzTp9nIR/fdH3l646OSry3dq3aTgT4G
FQn5YL9KCf8bnGZWP21IVLQHzCz7+6Pgqxn98Z6HCqZZOwSjFwctYm09C3TNcyq/aZwKC9jODR5P
weNsIEkhnektgjO2F+WOP+SCPwMYaiJO0y4r29Whd51V3QTFTUkdYsMPjAdAeXw2pZfYn/dVlVB1
N+co5zOMlmW0F4fQ0PfaI9FMYDot9A1jH/CHB0SPRUEC52qN+zYtHxXoKDlfETTDBvGnwqsZ6qmV
HV+kXgkbo9jSe/cGhCY6qmGe5NzWSmtIyCGpC1KlowJB/nnegzP2t1pAs3XaGVNgDhoDIFZl82FT
capHALFkMWL1KZ8lZl9NqWNVZLS3XqBbYgOIhAeB+ZS4yTtqbubH4LbRAZSrMH1g7iDi/AK21YaA
y/Xjq2v5CnBBDzCePX4sTQAVOaR5RQqHYAzZgrMymfBpXnRoA1EGYZSwiS6YdcToY6wliJXT408z
ZmCxXf7Oc+w9FvOp4Eap0zR6/M85QxBAWQOegtx3F6+ItGySSpaSzrSMN3H+pMHiff65psPYDtN7
oiulqgaQo9bqGL+q8RQvfvNLpSrY3j87D3dq8BblKTrf0FlMjyZ6G1ZBkM9feU1LWpvieNTjyOgF
Tg3EWi9jaGQoxOnkXV4ruFDH1B/q+EGpnXSi+0uVlPIQiZSvhlzDDHPPAOnINm5gNlLoB0b1Kvkx
A3rdLrYbYyyur33eH7ZykYFcTK5BR+DU+zgN+55Z8glocY2l+DRTalLkec1Rag5o/FoH5tI1Vju6
GDD8HAkNY32nNuXUfpU/93kfQpQtMvtAa9yOumeLew24c8/UFsRuWfZryZBJjjTk5hRpiuBwqaHi
cpSnVPMErbod6QL2YaaYLf4CQ1wciqFhc7TIa8GFSPfj8OPSS7TM4acSV4CjS2E1dYxg8ER8LALG
MvYzdmcRYZ4RYDFpeJ7BuHBUYXoNf2zG7eqWa3Z4aZyn8WTQ3rY067qbLUuhqFuYRkeEg/ddRICm
iCzvhVwL3H++GHe/ysc6Q53/uvzgWTmUu3TOAwFpFnUMV6kccgcJiiZO/vZJQA5fmvRy31mdTf6W
zyr4M99ThYsGpwo2ZmLkqw2R0L5TII6Sa49+EvTwWdXotTSWVVDnI/F0gVrSRx7wqYrVB6lpi1S1
h2tDt9WCzp68mRQA42oQtPviwu00cqpULmjbp4aAT3I6lOxOvI21N7LeJiDibeUQVn1PIbfhIARZ
DMpEkq6I3FrjuKSTf0qqJ3I+AdQU+/cRB62t4UDIZj1lMAabb/dIW7L8nnJ7PG+lOI7fWJJwJ3u4
zRZ2c8DTxXBp7AI8u30PVq5HF7VDqtlTo5WjZshJe72Gv/k9zuznHlSq1O/XH5jgAcRddsZrOGF3
SlqWOagjRWec7O+7ux3TR7dH3q1rDhcJwNf52k+nboziomBduI1pkmNOh67PLo9+YA7r50h+FUdy
wG3Gf5yxRvMnSrTGuDHXt4+HrWUfcrFhGJAXzN06slTm9OujCj/ntk9RTH7ybLecxbNXVHX8wE96
9QObJyyQt5twW+3iitWuu9q9qjGLZ06gmvbeCJ7YUpmDdzyAgR+YH3mG977HiAPC3bYVYlALM+/O
2TqskcL2OB8g+DaQJstOqfWhmPGZB8v5WNe0dVDk7cg5i69Oj7e7EeE15z8ljwy5seYxTmkYzO5K
wUr4Img8WpPcu4stQixjVBHdQNfKVwCdxb8Bsal45PPd3vzmrFQrOpqFvoq3g2gsgJRiSxVEUbuJ
XE9zlis+WV6FmPm4S/Roct9XqQewPG54c7mjFXd0kSj+sfHuUb/zEST2epq9BkkY6vGV3unmwEKu
pigIvYhguO400A/+NdmXqekiLLLCj3swn1+aVakLS8Ox3/np0e+9PBKrm1Po+qm80T+HhnyK8POs
qPYKSIi0J77m922KPjDXanGAUPiSHXl0njoOq9+gsq+kbVFI1oSaj6fCHUGMSavVoYVB7CdcTTSR
0pzoCJGol4auKrE2diXoMvbQSW0uL/kuPwRBX2SY5ccLCDc7l3He9rVdEEWF6XlO+LxpBt57ZhLT
ZYOwNLW2twptNT5X72kzDDx4qzwF5hNj5ATkDuP+6PWrow7ogHVcOHKUYCRlbQYwNYhdw/bUzEhu
1jtn50/xYCl7OPWV6mmbG51y/WMB93yoEleU4OnMDi5p/3V6C8jJVaN33OilTTZHGkZaWVdWzUbQ
JTURXgQZvklqfqWRq+sgtJiP1q7aquUAiqLxYqg33a6MXWqNNNKvyantJ0/XquqrfZcfIC16mn7z
SaH+pa37wl6e8092i/sUPtgvsQdN2SU97AuUyxfsaTnUW9dPI/LSOA+wWirJ1KEFJ/m3q4QB43Z7
JwYBvjlLgNPvxDwStmPcMZnUzKFxp0yW2hB5/cuqxt4WlNGSkCxyM2vxsnAt6F9IVVVB8/8zokaG
AxaiRetpCBMRfUa9CwHqHSL+bOOLPmmueD7KKGKguNlaCN+IUK97TWGmgrkWe1N4t8vecsfJPkn8
n8iLVoyzGYcdZCAyECmGwAl8hk8c2LC6vvqcZk/J/2YK36+0Th1vshzjS5oHZovl31PC9xtucGSm
3JekYBrWdtNgnVtnF8zpPalh3/DQ1AufQ1Kcdj0skv7Kb0bSiujkOSc67EtxHmzUg6fJthDZHN0I
jdR8r15ik+msj1ZOSRwtO2SX+ixD0sR90IbdNUhMVd4zA2Qgl8d0gQbIRZRGjneDR4P7qvLSIyyu
lFDsPCTxS27MnUBRK41fGwCr/uIefqPXe5+vx/ZIVxK+FvqMeG6qVH5xOTe76b0j7be/nA9lNjKP
JJv/YUMOZ6c1R1N2pPs/j19UqSiHhcb8DEBi49fRDkJ2m+feAwcZJHW6G3L+v44H1xcX5BzffOL5
xK6yEHYx5uXobB4VPQNelv1MyS93Gv2Zh/Fj2WPONtFkk3Hvm3ukIAcAWuHt3CzLPkSSJ46TIXXJ
4Dvc+pxDt52EG0gl5VBsgx6zkOTd+4CTuR6zHF12X8JyiAI9Axr+H8jLCA7bp63lDIWwR/nyGo5k
WLpBYpQ24BBkuQ+KQKDsDK7Pr5loUO3N50SZJhE0XugRghtZ+cArTrAsWeuFvJa0//LT2DKqUCCC
zdrgxUSE2UPz1ixJN13rPBqytn2OlwJFHkGlCDfRpaqLnvnuQhPSTBYwAoQydu3H7pt3fadTTVdi
LPli5XRVX5CXplkCauUlaKj8YHwgirAkwWOtSbQk/oOdMGtDHbfvyx0OT1F3hHz4dds7SnShC3u9
PmWAAYGZag4T7qCSaoRfwAG4Nqvj18CvQ2/xT1X3ACFyVeqQ5hBy5BX/Yv4eEkwIXp9QEZQXwh+1
TUI9wdnh7kQoZb6tvmnh7M2An27D2nXbgdJED4Itb6EQzcJyjkAYB003HoY6LwNGyuG/hosk+IPt
ddM22X0Ty/GhqZ0nytuJjD1NKoAJkJHiYIGx1iRbMeoAGjODzxOgaiLN16d6lFjiG1SVVosb+xwj
t48Hd7YDIAwqDSrt8Fv8Qtk7EKBQctVbvi5UB3n2jQjwELkrxDc0UfwDJSF0dHqlzPasbIzMnhiq
NMcF8rTXFM6jI2tzWlZTI+cnP7ZnsjWDL5FHwWPTLGjtaXmb91X5HaOnVBktdXcL/Np6d2qkSlU/
DMCRBi1RY5EMa/RdBfn0yOuujCdbsk+RswR7SBMoQ0PDzNOdunA2lWPRuNtfd8RVXfYVPSpqwJNv
+/kEK/fp340CBVF02W6c2bPVjxAgM03MunxJTRECbHSFi57jSWjNwXbQb8gBkkGxVxQfUZuB19kL
SdZ+1cP2BQQxWnCw23u6pq6hy930vcjCHikMqW1lmLEi2TlAUcn6mkrVz6w1KIJehIBpIXUbUiNW
PRj5rm8V4yNGzh9M52woTlBZ/Y0n2WJ1EwyDwKt8SpFDad5cZrxPYIdpxWDAmYMUsXMwFSX8uEXj
S+zWG1FAdt7IY+RUUJJ2AheFv+EqrewvmIR1vF1P3FFnSB8Pit6y2mVOJ4E6asYS2ZV5PhI7S4PT
ywupjprhO2zo3/kr/HMV3BXTeaVIs5CzM+pBUKZ+xs2/oBPdwzobrfqplgLB3BnWtcXXMte/Rcne
huyzOf0KRP602lMZMCBBlSeye6NnjW8gejrA+WymFZUjKKiUJ/YaiBuRpk3ofMGmFOS2dBOCqhjc
oYZNFDIGmLDt7o01YMpgFRpKdKIGUEqFWnP5JZUrEdtkw2Zr041NHdS0CkAzweVgIUUmeiE9v9sE
mcjVsmZp69xXQYXOJSYZUU4LT071wqPns1C3FBLcGuhp1PfjQcFISASsO3Rbqic+9lTb02r/+I20
0G2IoIS8ESuH5jMDpGK/4iUnjrpB/jUkgqcOs4WYoM/LrQhNh/Itk98FVoOsABsGOxNIyK4VcCq+
ueztP3W1br0Xpdkpk3GgaNiFrkGB0nYIvlfe8xz58r95bKArPpd4kG3j7skNbGn1vE9ot4geDnCk
bDrC+RAwHbT5LMPATzdaCGt1vrsN/lklMkR2Fht4qkFkW9EbytfT+XqUWb8kOGApRciYVFN/lLrQ
8Dgr5yg3sYrGtL0dUhcPP+5S1kopZTV4cyCaksDdARro/ax+57iQIZ1dLeN+4BjW027sIv0BxnvH
SbOv6q/2TaBBAbqa1ocalweu0yVNg/qSYypP2H3ZOD7lsnt7ViFs6QyAjeIIixvJAKU44m50wB4+
4v0VAW+Qwf3mVeru2N+NuX0MRHbTtaeQdY/YtddlH1IZw6OT1z2dSphZJuYgNzGFHSaMs4THiw4O
p1Y12786AFHpfrvGLqQi1Ic8I0J2Q6W4FoGERJ4h4FZdfx4YI+eAVP+EJH1OZl3o1o0KIjKy5Q2W
CS+HhwPD6DTlDPHJhZ6sST0Kg9A755OAuv7EiJP01ukVzNrvdEGpEmg7OriaBLryM5x2DqrR+KPX
qZebfr74qIklLCaDXXfZhaZbfDfnmEbdb3PnRKR00O+US97qm5kjsJqk15CjGxXNpMRt5N50ULdG
4sWDynojyv6O7hbclMHBdX2YmrF+S4BNTb5w6fBh6kDaU+/B/xaqNpxHnk5kM0I7uwsn8M6pziGX
JKTuKjSzvUlpM6QpUs+EJMikzXPR/aN8osumuvFLmAXdYPxFJYfvc4jjtPGCeEGjoH4emOCpqBfo
Sd29DvBCC/Me4ARNFh+3GM2I9ba9PUVRDhfZKheH/dFHZPVjPZMrGLm2uThQdcRHB2e1jTMlESLO
G0JfFmqOF8oNwGfG4pWBGHL8PGzILS265gJXSaqCnOyL1mdYrFa4T3JsnssMnLHzRtxjEO/Sn1vk
9fyue0+xgxY6cgeui2XukWwuHp8YzYhNQ0f9akIwtfW7KYCOyTIxaKxaaJWr9RRTw/pP0mkBQkG3
cCZHxkwAoWONhDS9z7N7E6MVtiwBxW83kjqtCM2JtSeJTE/rrVG3lS7O5Nipuz538ia8u6/Feh8F
huyORCB+wdJYisDw99owmYWmnOiloev7o/zzW0UcfGZUzJ8iZr3HCyCZMItEKNByK2oy3XfdpSQF
DBEZCoFqsTRbjfZwfd8g24+VmsKU4y/qfbVWRawnNv7XnirfjH6Q6NJB29yoMsvtyCe8+ICdEiWz
sEeIs9jGWrvXrSglI+1OfHCh3voe9Qm/MxXXo/mnRDLZ1OPNiARRBVNJ+4+KENPAZG7pOJa6a4qG
TgN4KXB6z+z+3V05xpmX7ZRiDbvo8BCwND6Ovu3eakY7bcw7M1qx2EZ+VUVS8R8C608R/eKPZa2U
PJ/tNoAvoIFDaRE2pchEY5cnIfTsCJysGL+YHlHeM//UvsYXFzY4KfOSQgoYgMMbM8udCBMvO3Yg
Ii6YvU7YWZqk5pQPipNJY70hdpGJmUX5dcpfBxgDkQg4yE6TjGvCroWIAl/Ytc1y2YelFskmfmKc
k74XMJYQ3myIVkHq29jkjt6UnJEpcVEVTFDzogqfcXteUOY7Vc27AIMPSkWZjQZk0/FFHXZKYyx1
lh3ZbFLvGbvKfchn8APQId5luRQFsmdt4w6FozbJUw3l5UdPxzrH9+8zu7yXYYxLzR/iw4w2RkmR
nOfBrRevNJKAjqWe9L8x6cREBJsjGdVO4tPVduQPE92qJseUSaGMP24HVMS7zUVIWNueMD++DXLj
aiF7t1VJAWAzysA88lK1GL/7V9BVsncTQDSNP3SvS4XVdgBH0BTSLoSyugzXuExKEKPAIcsHNSxP
dZzSQmYIz7T70QsA+zrMPpGEmm1yBsgF4LPinU88phzb2ogcyMoLdk90wuVudp+cvmF/eJwHaetB
/OQ6FWh7QGkll7IMHPXPHhJCPaGTfgrV671bcEb8e2XMUtM/ZLA8vi03wwN1Lt5j8mYHYj6OMhia
lixTIiz1IVRtxxDho2Gs5cBaWaCObp0SyCyG10AMBUWIHFYCNTAmI8lpwM2qgzRKaA2/9rqlEvU+
RoaBYKeFXUE+W1D49VHY7I8UC2FXLg9L29Gw+XXOdULW3PTs3T6j9cSY7f0INNwcwCjBSNTKavpb
9sUjsF9HBugPFMCeyjQoQmgfuxbDBTHA3FYRzqlMx0HobggQYns8i8pK0/13/UV/gJx4YOwoovyc
dANJJ/wCufp/Z1cqwgy8i7aG602hyd5STo+tsqp9l4J6KxJDSXnrK81s89xxK5PFq4gf7o5uz9MT
HcuSoFE/S8SpYZC+ssoYJkR7K3cuVpRl7axOfnx27pPbYy5ehJtPxfoOnFdbXw0af/FinwR0hZJw
w3JxgH7j/uD4cqLmlMUY+Ao+65LA7nMqOBVctKSgsqVAgV2j+wTmlT2bSPdcFfSnp27I/anysAwV
IiPZ2GwilCY0WY9+1CB4eHA7SvCJEq4Uu00pXTfd4SMrb/HGr1VLWRQQKsxisTf1aZuwg2Z5o5SI
MJ+7QQAWXMNcJ9MhR5xtIz0UXNJJJCrS6R8i1ZuvekIHZJnUnTMIe+KtPEyaqtv3vScGvk6bviLD
fGd/uFSIRN6D1d3+Mahyx2dftUrHXfyx1TSPinTkL7PFqzBIuX72syCOyoB1EJh6+/lkv1sg6Tix
7rp/6CfzNC0VS736fXhzou+wOUW+z/88Q5vNKvRxpBGrCVGkad9UVPJ6NR01asl7UF3zM2tKW7KP
BwpHJV9R4ikipJvZlEr2thV5zmggpVSPSopTVCqKlnRjWQUvhAenr5E5FG5nUyG2GOBRJQjZVD1B
eGc0g0rCVtm8MeQQLhbgrc02/qht+FvIUemj2qUkZceTVVxEF+Tgy7HwWoRveTDlwZxt1cGgokj8
u0i79TAVWLQx+vkM/yGHgg4ZeiPnii87qLSw0hKYlNc5UoLj1rFZuqOEKITIC0Jeu4kB9M3FTbbu
DgUR7Q8skJXNAWxiVCFF0LYbc2c/N+rRfzmx3NHw0XZYBciz8TBAx1xAmqbcYEKpRlS5VnxY6TyL
UrEe5/tPSyNJDc35c5VbKUR7m0EVth1rrSp2u6VRK0z0AoiyxF3bv+AQuiHcRIeGlNlboa5AyOhT
VDf2fzoz+yGohIsPCgpsELUiIkFGdxQftM2XfCbKxBBcIxHjjOLevuMi01y/7XFyKSb89bHq+cVS
1Vu0Rwo17lkd/UBmSg+L/RJUtKrgHIG4+YkxNNhg51qGIn7avKcTYFtu0XqzPG4Mnxi/IlDCxvzw
MQ63FOc2Mz0JjXHufBEOZKaInNN8Ahdcrv18j2uj/IYmUEcNYLXWsrBIE6Dfkit8Gy6mHtkdh33U
ECUBd++PrLx03zmrkpo4aCtVy3QLn0+dPN/NFJnv6re7pCRg+h991HG6jKLbh+H/oa6qiwj4f0cQ
lWUu0M9XlfL99iQVaRfk/WsqD3gwO0Em6mG7tw1yMj0/xg5QdVkRnZNreH/P5UcmPTyxK/2XBsJf
H0llWywQiCofyAY0UEX3Sy5OIFaxgSg9RwfKKDVpGOmwDOcu+/oDdVRMqXVvP3nt+EehIJnEyEc0
2qbTwUNKt/cSKlr3+beF/DssLGBtXDfDSNHQUxMs37XjOtuKVxffBFDNyuI7UfgHUlrDmm3WtnTS
Ff6giowYUYNaBdj2uANf2fUnIy3tMWl7BgjLUhOxlnmYJZUuJK0MgEL+XzVI2NHjWKyohilO7+8n
CpyV8uz+OesA/MVaBzUdrYLpJQz1chO1qtqquvzVDucI5vt1NYsz7Z3p5LKTYc3Q8/QqTSUNDDhk
3PRWnCpMLCY4jNsdJFSTpKZNyS1yOfMMAhmgTXWGnicFsxbJ2wEUhUFJwwX85HFm3cYs7yWwLEPi
7Dq5hf1GBSWlZokDI+E+obI1OAPuP2s7Nyt4rJ6uBnBir0O4Hvw3SKi+Sf5gHloA8R2jTri7HEQD
DrPMBfDgXzHIiA43uLgN9/UnPKXdFDzNHI1euzjufBNyBL0B/gemDw2gu+lAoGNS31V2afHy1aIG
39+yTevsbrkN0IeBAP4X/WQ8fqp0UIzdRfe0BDFqwy4SHXUvCacqJvaBi51RsC6lZ4sph16zG24D
0Q9yD5odatEJe978Gqv3h7fbuM4qfjXV+gtaN8GBycZrecbx7fCIIE5j3AZedZF+RghVoU8q5GgJ
wj7rXobSUC1xQM8CPTjEHEfQNorbdrAWawww7tTm8J8/jWFkmeA3NGg2CYQOhPcN8iHd1ozLqeTx
x9LgrRnEWz35f8+Rmj6mzI67hCNHgehBb5FQ41AORE3Xel5sQUJMoZh9LkTMGGKBezrCpbfHwV9z
JL8JH0+ew/jEXqeb1+vcc6CBcb327rFNqs0HlEPAloyUP7LaA29U9JZ1TLMMDAV6QH550EfzDSLg
NzvSm73dDQVWPKmR9DMu3n+1kHMs5U5nymjafxRbaHRFmfLiZ2G4u6VjFLYXzVXGbQOu1wzjgpO5
N/+BhbLmWaO68CvBpCqWOB1cHdQWIz8wuqeuaMygwbtHSsMWVj69LvDy3Q38pQ4O5tV0BcA+P+JU
wVJjKj41JhoBzgxHe51WZGsvzFDbms8PPObv9ygM1x78OeKBwn++jSbVXmkHakmbOr4cBpnBHhxG
0J57J+wAHK5Jx/RNDPn7KcYa5RS/ws444oUiIr3boSrpCGtgm7dENFY2K8BzClq7DdlwVCuwNq2X
y6r+oWwji1mMegjzp8fVso2tVJl0h4MHqFmqow02bQ8Fy2QsJGOOCMLxA+HKt0n4NE6E3j0libYw
3LyI3+VOPh5asptvjLvvSDq53a+4QXHhZp9+l2rCbEevCHXEylNlkHEvlNtU+Jj+myQMAywDFx+R
eEvAwYKbUoB4fOGBBxw+DKJz+C5XqbOfD2Iwf4pXkitV82B1LqrB/3u511w5J8cZX6P3T3sPAeYY
ba3XPwa2z8HpIwrvHV8rBXvHmINlluUejPcCL0NVvYlDYGe1gjoPBs/nRf28zXbzXa4lqwiGgUzy
BSTbB2b45WViCrj7wFbDmIxxiHzhFjsvfh9i634hlCuH5gyFpgMIDv87iYsnOgsltxP7FQOcju2T
0UsUpR+3t2IdTcDLIvXVB6X30uMc4/e8khi1uSUF/PFPAsEyUYfIfMBCYw+ITLEcGoHVndKrLfHx
Dx/B7NpnEMOOhTZpddXsEPEXnTeIh114A96XAF87LDFABrVjw+uVz8+drVhzf8GyHTf7KSl+6tLv
FesohVAurmM5iZHxnhGml1qFholck/FxA4Kbch/qS+h3kOjNlFH+i3rcSCnrkJ0UHT4AJfnFLnY/
WsoPG0vVdcZc+pO8UGGqDF8CYhtbbQ+yashSFx+CC983CscdewEqjrd9xm+ZCgL+yMV+zn+poiwA
3tGnDCrMSEriHnneUW1Y16tpMSVk+h+qOV78op+5g9VSL/gp04+KTHW5bJFFdbp7/iGp9QE1xr2y
OVWkE5rP+tMB15thKr62grNtsWPziN2aP9YfgF+NanpA5CAX5B/cn/eQQvcoLXQ63ldQ52CLzqml
jpIKG75JDmVYhwdwni9lPyjRHjA8jFJxptzku/d2mRtvBfVvuRqISUEJ/OQtXtA1d4OpGro8+aMv
8DM6cWnPIQgsCoZ+dJ+edn5hJBvUT9+2ab9lccmL/xlXOvAkLmqA9sf3O9tkYyhGlO+l7Dheo5dW
eAuRR3qBEpeo3ZyuGTF45Fpbn0F/W19VSJCEMKUTqdM+hOShyEO5lyA6tmopnTaoklsXxBhK1tKk
kd8D7BaXYY+LtRN0Xd0Ew5bSdIIDrvetQOJ9qVGaFcIyqD/xa9dXKeRm/4ekiVQ3ZgNW/KSiQL3l
ZR/agbUM40q6gJrRC9iY6rXowUv1vGACWidUlz/BxpSp5K2irc3/LIRRANMbv3VS1zQj7fg3MOEr
I3/19pbDmanFgQUepIjU9VVVZ7jU5QyXm2VXtzsCLx9ENw57WWj4ACSQoehihFxkch2ngbKeYm/T
JkWj6BwT3J52Nl0ckk+3o/9OKFMZ2R7FAigsXueK/lDeeTrek5yH90aXd0bFSxWwJveyfYUFAqmv
8qMSKl5jmd8HrQfdJY7xLtVJUVIi1yIothIpUe8SBq33Jj00EJEPpDqr16Wl68sk7n7t8Wzoal5W
C9RpwkI0MRn4jH2hKpxnhE2SC/WRnvrt9NqrJCiN4L87bR4eeARpssMvRjkSMK4jpMDj8OGea2FO
/soqnAwAfuN4+ivcXJ5NopUAQ8xZdTuLwsjEZL7yd7GEIK3R0zaU0aGygVty2vql85ofLQjFvIZu
ckGRlgDucjQvxc8+y539tyBBCXTnOJafJ7nqFjBSD5cLqDoSJq68ut/EtfCymgjO4AR2MA/lmpqR
xHMz8kDS8camD5yvnwm/HC1e6I4HBWK2d69oKdkP2gbPWdGPxG9fqoINDEA+mg9GzOj/Me2oanF7
1hv58ZQSuqNUXEGlvhAYn1iaVQK3zfymP0hKyoHss3k2h7SL3LQBYpMUxhKD9E9xJrCtvdtTHWKa
HKfpS00LG1lJyav2Wqgc+fAy5imw/WQcIGFtpCu9uU4pg2DcpRczmQhb6kzGcfp3jd32Qe4lNa13
Ax3RSZBvxj2e/D2trlUFnU7GDnwZ3vTmaCx1zWi2hbNDEfow6AqPcWnPEHEN+r/fLFRPf3b8Ukog
8CSaz/u9TQ/ceCt4WC0WLeRq9Y4xSNnRalqqQRXJe07L138EBydKeX0kiYBUNWhX2QPE/gknd5Z7
y44Y9kQlpKUuW1g6eVFhrWO71JwF9EvRpOmE2H41hs6UP3KvMxHcyvOlwc0PjnfDA5JFTCGyKgQj
eHJGOTK0MWWb5b2oIhfZ+1ra43V59T/5yIxaQxyRCdKiZKCdR3+RHQzk/bVLmwZmfXHGuF8JPmBS
qlLOcBWhzkvjF81r3bkajMkUJVgOMS9ylkGWvGdKAyARIfXQHTm+VeY70xJzTdDcSrvN1ffez41l
7pK++/w68VF+F8W8SGFRwxX+hKmiqXTbJSQWtwNvQO+Z1rHC3UzKHBoHNvDEEXlO9Hm3h4eDjZ7S
jtacNdfn++VoiiWombVuMcM9pPReu/+32WSmsXrBg023X/3LsB93pt2TI6PtJ2dKqujaGekM9RlY
SV23Jt0+iF02+Ept21PAmALOlGuKvxORCSjuJs9P4bBbOlpe9QZQKKj6OmfFKwIGPacT0jLNkHrj
qDGfYEjUD+IUkvtKSm9WRNlYOBk6yTrex3QQdeCMTESWEDatFXjlQR+tfCUJJ6Vwc0DIRH57xGzS
99CdUgoNcvTD0j3sivSd1Np4W+3gyUA8/EzH6UGvIs7uQpH5jqBtvTV2hKBgbIyGlQi3jNlbNXMu
1IuCgl2yZM6/U9gXV6tlDD84h46qCLJQP6rTtaOmxsoMRWjdevRl4quw9wjnx/eHoTyPZUPYmdBc
kMkX+CaVpAxXFZ5SFnLiVWBMN9Qdm5dkP+aYUIn9pnGnGM5jqSWKWAkuFMuhdR2HdbGKYcYoaH1h
6f2fHbFn24K/cKgl7aUSNL2OX2sxlrASNrI5sUF0tUoG2Rp5HI2rUQH/9psujCPfXf6r/tWlVCYZ
1BqBNGKDE0yDti5ykqMnaETaJStW3KyNizUszj3M4UvrWRPHpEqPejP3GgfRj8k/Qiq/GQWiujx6
YVgJPtidvXy7W2bAKshlAsCwwbn3SEB6arsBx8RQE7mONu9PVDoUMRt8RfwSzU2WdLHKAsVuHNOv
UvZ1+ADGdlGTKDc8jEpAhQl/i0/mrw68sRTjpLmV1gA/qZUOwzIpcLssg7+pYZIvXpDW5OtHekMD
30T7OpCX76bDVLxrr1z267gdAjs23DMGLSitc0R6cS0lGCXWVsc7ddtCE378Sw1hddOgRfFN+SBE
7e05ecO9Uv8NspCypT8sTUTIrdeYeCChnZfTWF/08xiV0QV+OHonQjeAlyNCNLchlQxIlGyDBcYy
w5A0FlR/k1VNmNO+Yao+lupw/Yi+BdtQGENzcfzaetChhjram0ROhLHYClArSWbbm4pcjC4Ile6e
fZnYo5ZBRm+v2lRoGUn9X6/5N3EY9H6NqUWV613VK/Tm2zTlewgUedmS2y4be2QwipVDrdKWWLaa
Xh/6qCBzKQNPh2XZYqAmAsXroWBCHfImGG5gEizUmqAacD54RIFxYjZw1kV0OtI3+t0dqfNsZzGP
Effq/TweHTsp+jAci4+aAzNnl+EfFLp+EuUjCVugeGH/8ZT8xy74QQbu4iZiUGf6F9Dgtmc+Fmi/
N+2Cm6zniWtMi5+B2l9oW5upL2WiG3tp44kCefbosqW/72FqdAX6RPS6uF2bn5J1OvmvE3tKN+eB
Pj+yYaO5Q3R8fy18Dk0trljB6FKhtByIMS4kXuj/Jj7q8DIFgd8OR5JsT59v8QMm5Goy/G2sG+js
EHOzgQJfvln9V4dqY3vB0D4awFVvic36du4Oap273zgJJFj033d+6XbrFrsbXnMuykPy0sMoh1tF
4QA2M25W3oOYivn8Ve/qXGeHmPWH+d5AMhMiYwmTjKXe7VAeBnJUNlc3PP2A+zqOqw8X0Mp3Dhtt
M+yThTCwIOsiG96/sib+1AzlhatTZEIb0o0SpEuXtawsRk+epRzFk0aSUBW8bZvUcBRIwFoRmy4C
johQHT1fWg67mNCEsi05NgCSVzhKEWWqUbFJLrG4UXRZo9UBEvjNlzWQczqrVw86v3PpsCD113aL
W66O0vNpm5sBAyHMLoLsVv3KSPIgCDPT57pHdijhqnpK9B9eWlZ0M3E4yVRKDoDF41HWtVO2tCUm
GteJlQy1y6XHn3d7dgtwaxYeB0oiGHFUNcITFUwSNfLMYj9soxb0SgZydvEUG8/U6ipAKsbh3Qjh
FckySlE0gbchzx2yT+OuwTo9BXYC2VJHUM+cOEl7BmYBDZQpJUy6vpqbQgGW/z1bxCTlTidEVmuM
44iGoZHv6eoLIVxm6OGmtYJdSyN2BpeVfDDjBCkR1SRCPjgWZ4y9HuRf6aaGT4jMyj7rHfBxfvVI
p5v5pw8dBImRHi9HTxtzetaZduZn3HdpRPSxfK9RcmOzX3LPk2E5LmJHzSXvBwnaeo3vDk4H1Crp
tf8Gw0Fj9pEsvVYpwAh/1rADB5V3T8O69UvAJluEjfBzfl578iQOWs9veJMBP2WTddRYUcymcHB0
/xxy8donH0x5yz54Ml6ztT+oxHWOePhmaGSM2/MVW2S0jIMmgTZdXHB6v2tU8OLcpunb/YGO9h8/
KiZmVji+x0y9lsWKo/FDg82+e4oeWttJi7xzT7himJSev9IvEQcKSdvtwZVoz60Kim8pVuTg1mJ7
U9PZekJw0AV7/Iia/Q/9LmVrpRmI12JpOKWpgpIRJBGve1lqgfc+xMXSKgTuS9Gyzi00o2n3PVnd
be5qlSSMVHy1ZPlHQkw0MCshXDxMocwjpWnvf+A1Fbtk1pSoQ0MCuEep/rEUs1mBB2QrOlU1MD4G
WIcTbI4vFMq7QIzQSNpWFs2gpFvhWQIbigdb2AHgKvTa+eIice5d+8jt/iNeGbRCTATxsjkVfb6g
+QH4loVIF6b0djtvfhjMUHI6y/I/6PsmAa4LWt5ZeAEVhjdl1IoPfAyvgcA3jmhHhY+0Fkd0KKYr
741rhX6BPDWMBss0NwmjAtrdPld+a/Fk1VeJPgMrOU73ML2EhLlj9sdUK6HtY6ESzBtrCJAYgZwc
BiBDnwN/fuwHWiczah5HDTifSFq90TFEDm/eeo+BvDg2CJYbocCzeGmsk0vO+y0+fS8WXDzZmO2Q
kPXNGa3R/6CrCJX2Xc0LM+qoPuXI2v3rnE6xT1hngU+D0H1u2RqY19HQCdeXHsbvnSZ0EQgJ1y05
Vc0U1/JjhSan1ZFOJiPUYcHY/toXuTz5MWhmQKw60WLeOjDkCT6kHDbvwrUxlm1xU/ss61HuSCRm
hU1eJs8OtMDPjCWaO/WweR951JLhxhq2gx0zfgEQX5HNddPC4t/h24U7EddW9pLF3MtW5HWCols5
qiVqgTZb6QtwZLp4JNJkd2qYfT7M8uiE7JFIA/Nq4MHB3KESrqh9bA9+MtckB4FgXDr40CPUQqhb
F6IloQbY4OBWCiMNeN79DWUxzY/6KiCwDzXkW5OwEr8Kuc0qZQZUsQFb0+aHMnXRYzS3bcOVJKgH
LxdmxRwABk7N4aG5I8vYeKg3zRJX8o0Lt4+vXvgdYacBpTcfrCIpzlXQP+eH1ZYJFRz/rvZ6H6YN
EJrjebtstOCUt0SHQDpW09bDmckF+85bwTd8j5JsfbhUBkNwvUACN1JoJoiMZd0dHUJgxsy/FRKp
te/VbhH7nQlyIEiqAUvZ3nIYB/Z56j5ko2bfjA4M/pDQEY+3bYfXyRjChu5VJ44LH68AkE/tBrNH
nAAGSCDIiHOw9nYRqwD/NNcG47W1WOFJLbfml8uQqj7on4lGlGz1ZJE3LMhTWSPBIuuuij8MinDr
PbIIUNq0cXDKY/NFRD2mIRlTgP4ibX51iaS2hoAQNSX+tzy/a1SxWeNEUXH7h3c4+MM1zQr6Xoc+
FWFkmSceFwo3Gag+IrhVQNrSCMRRmXYL6ym36c5yLhTNo8e0rHvvTew6bKi2RhZ/ymfArb7+V9Ur
EoySVPnAa6HTu3uWjyvInGUc9oXMon7sCGGEH/K4wacU26nS0ij2hHLuNt9P1JVAXp17Tajg4T6V
y+1M+czXXoqVzeQVdtSDHki66iQfHDzx2eu5P+swegK/8CAOisHooA7SayPCzhmLytSqZ8gy+0YT
PWq591WLmw3xgxQR5qa48GxitbgNF6mkNMn4luV3eeok5x2zF+FHkzuU1tKD1JRi/GXSMNY3d5rG
DVs0/+lczozZhN14cQZ4R8JZh4ByYrrFK1GLqaPAKemgwnRePW326dIGE5aGERrf5oudIQYd2qSz
SusvRmVZKRaiwW7B6aUbdmipkypG2GZMHiuNNoPnlLJ382nfMq5mXEi2ynyy37XO+BFkwH+ET7rt
Ciu7CyYqYSldw6m0TuZOupmDqu1I77YahZzxEIQGKhDlA0q8XlDmC8uCc0YTai4tx70s6M0+8t+m
tG6vBkt3+0JK+BNuM4Fh0j72HENyQwOxJRTYoX/FiQvER3ohC3H3rsrwfqhPmDxiJ39/uLu/l3sb
9dITboQXpafOyTSFfvfr22JX8dDNJmPuF0cACv4J3PC96u03SHzWvgZxd9X7AAcN5g3iYVeoyUDm
qSJVjxyHbD3hM9mKnUoOgaGra0Mo4bSesAxcdv8nFevU9phuRCdfcLGhR1BvKcHi2VMt2M/yWmlc
r5U94jXc2xCT2zeXMtI9PK+LOdJBUj51IpJ/o7RNSI9ljJ2ICYN20N445J2Dai2AuQPfpKslkP/I
jsyF0Q+ztNU1ZC3ZptTZud6eCpZqy/0H8hb4MFunjjKA1zhp4w0rBOI7T4VUKcGQRAPfGp4oPmU6
XMyTmxN/yZPCIcgWzXfVn9xLOXZPfvtlF/bOqCsumyFyWZCF8kTp9ZETZM/jvP0HeNI07hpKl6wl
soSow/SimeiK4Y5Oyta9lalIaCoGMt8O4HCBBzGvHQXTLeg/DeoDx/FbxHV3jVUbM+tHFCugEqVV
B+zQYRXAQiBiLPBP1I8hTSd07xzSQua8rCUPrOvv/+TAiqYPa6apIodudbPWDy36fMfr9llVrAzc
+v81ze1MEoTaisWEm/ScpqKw2TkpalrjSM64kO3SO2GhSYiQotwbX2CZXe7F1HBFIPEz1tP60FOU
iCFtSQq0Fo/jD8qcpf6F6BtZirTO+EKyprtSS/bNmdJnOTnMrgbpxysseJHV5M3gCd+bYTVWkiEi
zF/AdAS9QdpdNeipp/HUS7qIyEGITkxuTAPtK0ze4AR9Eu200SckrbORQQczp6RTBi8ix2Cryqrj
DhmJAhjoYT1J69dRN7mkUrnacb+r84IfGGH+OwdPspIYFlvonCCD5PdLKNkSw9IIvR9HAuK+MddV
mson0+tB80IeqmROeV6zQzps7vmTKWUpu5Rn359Wi8OXDW9AYw4CTgvADlJHqxL9sAJdqjs3qJki
TR0f8UUa2wuqST61YmkWdnenyV6M8e3kt6zR9dqRHgfA/XoyeKEPw/QBJDoumGdwhpMQWVKrKoFG
b6ZPhKybOEE2hHYBqhGJqQgrRi7dFSEZXT90pFyzbikphvZ28BKPmrDg1qBsRsl6nO8Rj0YOx0Cb
9BGyWzh0Sf2zoxAOgpnZV8kUJiIhsPF4Ed3FvWhwN+7ooRUf09vmEt68Ws7mne383+gzcGfzNOem
IPqIAWn+NGjyRtTcrErQEXsq1qihJ0YMjud1DFQx/A9Xg+5gtKHka4gNRgu1/YOuHNUEfK138tR1
lwMxF9UViSg8w8qNgjVpzwtbh3zlkgJPqvbCaxURgLIt3FP5Qv3b5ZDVqEjk2+K+lB197LKhsJ23
+d6Erc1+l0Ux6S4sIYmuKycxg4KnXQ2U7YiJDngezlt/5pBhx3i3/pcdf9nbPSlyIk67SgFb1u8J
I2oWIiI1fF14aJOZ0eSnuxms69cRT/jBOlhrL7RZ/er2b0NIISr0cr+F5SGs5n+mfU15UzR5fjBz
JuHiIobK56PvopD/YrfUS4uKNg4SOXref2PKEme1/tc/1ZYC43Bc2kUOVPvXzjeeF0BOPCfbDZvj
doKexi1obi3oLR83xWkbnbyqpRIiKEtnIE8mhwTqDv09UCfb5LZPc2QtTmYixe7IKD2xmrXpG4Hf
urHhD4Gt9ek1QCzzHXc+M1pYI4Eed7dp6yzyTgUYQ3JnOMV8clob3pXNfqE5b6r3CvjeJOwyRqUX
Fn6yL/snnk/f1CDit1WDnM0Pps7krAb65QhqPU1hmBd0xujwnC2yAtUHH9iF454FWNPdsJcOG7jd
tOn7Sw8VDybJRQTfAqp5xxFXyjkggm2MaA/WuNiHQKo4PUeyTWMMRLc1EuEBMkI2QaMjn6WFm/3f
XZONihJpPv1TdaJDCE3qJ40EP7LniNBPrlDPpClTFgltj/Ii24JoVOXQh41G0BaTc2uyUIC0TDfZ
/ubGp3uCSBx5lRxoNmqqh5u1aAz8DsDdhfZ+sfGKwvTj5OrGYAyy3wdG2htG6EQUcPOdkjxngsV6
8/vEaiQGGkXXM0TKlyM5gKtESULAx11lGjmNSOmhjffb75gXhQdA0oMgSkKSgqUW1yWPMHZr3kiL
AosxK2nA3IDgTvpeMok207QNS5hjcsF1XIPFi2ee2EKgVxVKEe9Gu5ObzJcBFReucR3dmZJCw2bG
QKpc6+s8jmMHHipCPpiRmaQBwU3pHpIHLs6S50XeHKn7n9bANhl/2wxOwWL8rzOtIOnc+d3vGfxQ
vVkUDXUHuGJK8GsaKxAuz/u1Pu6ZtXbrzd6fUR4SS5/NJ5gqQvES9B9jkOkHjXpwYESmxGA1RlPE
1ZwtUSvqb+BuCu15zbOq4Kre/XblqJGdWviw5R1bYK6Lmw69rpQV7i1HU6BGv25vkRFyMfGzXFsc
qPNzh4mNgSLuajbDdQvhomAAuCF0HBUxDD+y0fZ/rpzIe6d6+Yx2SEWKYQbXQ5PWp4cGmt4ABhyJ
3n7QWqLCk848s5+jUdcIErGxB6NKosME6qkOMFYj3rHw/dQK3E/IIC2L3Klkw+5/m7eB+iOvjKWB
yHl7Qu4Qt7i1A822J+LZ6DlC6Ky+tHzkkLEOXP1TaBFOtqFRsYdRLMK5+gqKq0ob8kxj5guiF4lc
tDhdVuzqHZcCVs3OB3zhWCStUPmFZx3fjkvV0fD5828u6TgICVEcpowgx2mG8xJQJDOxT1IhicTH
KnBHqZuTIvOlKc3BuRYRJ/EY//p6wrPBZTrz6dfPHOn0jUkqmJacSSZkkm9qvQPNnpf85kuKjcvW
yY1vp5/bI43wLLeHj5XfqK+2Se3QhhQjNUv9SHsHpX3j5ZskK1Qmy0MIC7JGM9e0As+ZglSNI94M
XXoW7dY09tHj8iJPAFiCdrNC1pKQ31acOiiH/Ubpzbqo1VoeOp4muWFgoeKBqinJS6hPnS+v94gB
2Hex1WMpkylLkQfZV1gSa+ZDk9q+2g6b813ZSWcEcPuzYbDs/LSNtGiPJXtolSQJMG3NT7bb/Z+r
n+CwoMiSCTEPQI+rKY7p7JdYxUbhIrrsZCsxHgi8e7Jpfc75KK3jiGbnax4RcIf8Upf+HZJyWSid
rJmjWY4P8gYsPVbRw4G/35hqUKBBayx8S+V+qNBB+JOCVsbbb2PBkMqPrWzMLWEQexgsw8bzrFfh
YkrfkcN6u2Tyn+xeyb/So/rXhbCnXOTjsGq4PuSh6VfxezZ43P/fB0YOvE/P8nNmwyJZ71n60e4Q
NTrMNC7jmWz+eLD8SM60hpvGmAjpsSspn+NlkM/wN2g0vqM1XiZhgxU/WrOs7KwcReJR6WsKahOI
Frtm2Qg4DupsYbNppby6zpldqgTRMZepB0sCtmkfoYNlu1vRGTbxr3D67+MKaTyX9TlKyON88NPd
3zpEoJQqavzDkzHs0LHTJUqit17UODK3+rSGdOU+TuuG0oYsj8ngUAI4WaQ3Nati55cGmNVLPwLi
RRSjID0Optgc0ynNUr4YMo2rlwVirg8aS6SVHgaljbsp/84wJv4gqot8lwLX4QixUYPxeh0o/VqS
IY4+fX0f/+ybIRAWNJW0u5TzaMwbkeZxB5dYTnOuYxfD6i69lYYVsSN9TE6K0jo3jh/+eMSnfAiO
QLtjn/KEK5ULl4w8Xkc49GFyhOV8fTVVzCfMLQdSxzto0vPMyo95ltoHdSJzOEOtXh52d1dOR7Ik
sZGXvrlFBsOoPlDpMJ2mYzM16UIzM/w2TZuA/8FO9jFZp+c50vJH/U4lc6buoKRrw2Wdnres8lSt
BPS9LbJFzyKT2g83rxtMpG/CF6++ZhpjYznEq/BkXxdAWFjufhZeJuxGF8RgtEaMZ+a/LrcwVtkn
XGtGVIZYu1KUwg6+ED62P9cHAybBqco4O3BvalIcM0nV9QY+EnmXA2+PuL3wTX9iLRG92wK1xzIe
BfggSyyHO3xoAFWVEWnYITCjSbb603RTmIW9wfSsisf73KdjlhrlHXL4ineU+YcSC/+hk2hM75RG
y4Rj8y+LbwxpnL/B1drWllCBhpq2De5Hv1fngEd3V3TFwBuZzvSvXKvBLHNFW7wM2sc90JtxVx6+
PJeI8tVrNJM25lpw/E/2Xqfmq0JTOKIghgso42jSihGe2xXTJivV32ImWeJTFvynlagRWswH5MYM
Y6z1mIf5ts1JcOFaObffMcIOErwGMrwSyuYvwFlZV0COCH7EFGeZ1j8A00zEEoN+qJfLlr2WwLjk
/fQGaTe4Nm5AQ6i/6dIYEZgboY3iiiS6qkEDnur61nOy/6Gqe9VTtsZkr4bqtaC5nxtWXnz3mgoP
chs3B43TXaoPRvEWpvOFYYjLaauSb4tjmZo5ufYsex7zQmrYNU1MCh6cKEfv+bjwWGuaJOvm5mC6
505xHj+gBJVjfB0JGy7hAVMWABh4n0oVM1E+Jrg+dmoqvXXm09h8deYkSISiWO/ZFkTHIi6plhbn
9nn9b+ORk/FE9tfgwf+BhGmOhLvbGpMQv03kCOsfmc2EGDJ5QnLcK8SBgOVa3tfYuVeoH7vAgd5I
fGBKAKqmaixmFHDOrSK6EYyoJk2sD+yFNH40zqrvnBhqThetT7AqswKViGy4SANF8ALat71mULYr
EazKfSyze4wCS3fyqsdIKlP/UIcEpxXe/bM739A9vwRMAIba5fAcO1Gyd4cGOYHNTKTlKUyW0xlE
+P+iywZ3n9WZ/vOzF82T80OMtADphoOZ33VZY3Nx3ru1NXLA/K72KySrVm9LZxWsZ+oUORsBkP8o
GIkNItKExw0iJRfSKImQiVeZFEVKWs65wxNZ5FCko9+Xg0FRREen4yrfQeDlLQmd1LLV4KwNneE0
0kgLFaDrnmIqdvOFXu5qO8MgzB9oxtpz6fFGi/qoX1d6wHJSMtXgzw5d5P6z4CtCIm9skpCGa7ti
5ul0X0MpQvzfMVKsKp/o0WqHHQJK0WIBWXA6MLy5advGgumMxF4abFKqANmXKuVxLDX9hk+ckCT4
Z/jbRRMDdjvA9piW4t/xHXZG8dbjJEBF4Ws0ERZsdH3oc/ZClPPqxLxOOJwmAKYinkVGGGNxcZPf
fS8oT30bJFCKhpAmfTFTb76MVUNFAlVLK16XPJ5YyaIw6kZuCz+jjEaj/4o+MYqhMCEjmKniDISq
XYmyJwujR/5sl3pOUecV/MMN+rR13+YIMySkxzY6IhHnN6eONGHKt19y8Xx4/L9/y9YVhByAYNc1
IjrsO67Ig75OMgAP6gkBc0Ftj3ay+dDhIyKJX7CKcWUxYU/1kUn+QSF8jlV2O7uSWEvZTRyOf3ed
Rj9ydAsTBjJ+TtaerbYvd0EmTEW/bQHlvA1FAWBtrQtb40HpDdYvlD2pHPlHmb+r9LZYDc406Vpg
HgIGuB1ZXR4KaWJyfevmUFIHaKnzAunh2eeOabTbOxHHnYRpfNg5feQ1OcEgCEIsyIQmfhWoz8Ox
pyvpnrhnX3MC2RXtHhOgYpzFbZGITCVCnqfAiRCHHQdtlbQ4q9rzgP8svuf1G3EeGc+R1WCfm32w
HaqND6nfLAdgnN9dYaKWXtuZ47bCBos7Fv1rxx6xDQS2QU8oWG6sSc8hiywuyVqCwW/a6gDGgpih
lxNFriwxgEqtDtZYF+kKL0bCYya/qBwtf4LolsVoa+a2p3r0z+nN/yKDNKkpCuSk+pOQaPIZIvsK
nFgdakJjmGo1XnIvVFCLOQrL8XS12CNAt62aIlXtsRbdwcnYKolTs4Ki9dKW+gN7bW1mPTjl98g6
Col7zowdmcoDGjtZPX/IoYhkk9en8V53uuJKxCNbiz+M0gJAVR86NZmWLkoDtHikxwRk9OL3752o
IijNbFXfm4uY10qxjDtYEN+SQihpbAHPIoBqz3RIkN/69YsnmtRGETrdtsn+98UDYVwqT8zvZ5As
MZcnDj8XW6vDnKB54ikTgUWKjyxVdlXlWuWYhz5mJjDy46XgfkvNVAsQEe6LwUwJIi0xmnYH/Odr
FhRWJ+X59LYETInzwOvG9MDO2BK4mVWjmNPGvAcQw0J9CIPNcnZzhS4E+xq6ds12T6inzV2GC1eV
rI4oE6tcyuZIZTTMj0nSEHQSTNiDaj/2S9f27MZU0HK8ZXCJoy7uCuMh2UM0+9/qaohBu9sRN8td
6X1rDfPjyTk5rWblj0Sel6yAer/8/bnbP+Wfu7tRnYMT3T/baetLtHAKmDCvZS5Fu8agH/wtv2FM
FydWl4KlHfj/DG7/umiwaY5EfaR3LSPNFz09l47WmD7myfLAHH+ppjo8gEqWH/XzdoyaLkEq699N
SpYbGgypcG7bIozkV/gk7YT0lTYYCuCy5GNwO2WBSworhkQmEbT3PcnAhvgNS7y6eogQQ7riMfN9
VxEXbzhDtpJOQQ543T+OnWFki8/JYMqTNjT9OgqmOl29A6K+R9tdL8he2JsXzMo4bzU8xYB10N9m
bTJhiJdmC3mPKsrP+V3jtxh8afN9NEYiVOzUp4yY76DhMO2lRqu6JHy6eiRKLN2yVKpAXktSwgh1
p5iGqAMpvATkX5yORt/AEnmqxjFRPFfGdz78IiSgEjQjaABeW5evUmRxmodrp7t7aVMHAQ9gFubu
ogxM3UesaMm2821Efnid8JWQ0/ygi32LxHCL6zTXXGSoCMqh4lBSLoj5/JHabHNgsDIFZcI+vtGj
JdNYU25RCkRyMg54iVlMP+7+v2pJHm2LT3fZwIaXYu7ZLokE2G9O5SI0vxxPYUDVcg02h3Ctg6dj
VgGmG/FaAj7TMjrT5giuIx1n2x61VxeT0xbvwt9klIRUOG6kBT1Hp1/Nyv1HWvFTFeIvkotJCwAv
1+N529kFNrtQ3prFnJW9XmRSxScGb9DJDCG07w4ab7So9l3xalS76eiuoCmZx+ZvNhRd5OLqhZPa
d7UlmP7xnPTjasLnXgXQjjURqRTf4SnWQFvNs2/neXQ++nFuXefLnr9DDk+x5+Zwh+2ylZ4BhQP8
60gTUbxhieLps2VQvRWsCwfPMFGK/Cg0Xhhh+gHoOnkJDX7lzfPZIsMzCPxmL8LmXot4Kz8MppPB
mLfIgZNVMNvqvSnHsprEncXbG9j7Ho5ZuZIcNq1T3Joa/rvvWGwamD35EUgPRqAn8T/E4dEZGs3K
OnxZUdwRO/ORaeHxxdgVPBLwrHDhjUtrd4dRr7XiIBEO/5GM55PtkoNP/J0Gm3SdBGdtYTgCs+5v
e3l4Yu0Irg6QwLCuWmDOdE7eoMKI8MSKdGUGUZ89wiEdDqdd/rlcCbci7h8zKSrFHUU6vbhYd0LO
qadhQltHXxeOuPcNcnKqZMuY8uZIDLYiso177c0Tv1KKQSwcnb212OadMUrlUf7LcGAqcl55ov7u
lIaXgCeeT6V1klv9t04oFkDLiXkzgUXWc9PnrEQfWxYo2GrdAztHbxmRVKpxfedaRtElSy9VLNdQ
brXwVpMUWDxN0YtWW0SI+zMCiArHXtKQJWj/mss7LBKRlJXe7moRZOsvOiBqkfaitFwAP8FgOBlT
xgAjlBksSuaC8Ts7xpasyE4R5pJ5qftY/phW2HKGOFIKeCjQvQt4yWYh5vzrcqg9aK6myDeHJlCD
F94UHkYpap0GsQpBLM6xTWAk9nQDOywoY+LnWjIcqySOvCb/AZmrum8nn1slakeDfK0xhXxEpfVq
/X5cozVjSyOF6u3PjQaKRadZVg/+CsMmq6+p840cO8Je4xQbVFL+KLGQj1JRLAseslLbbq9tbo5M
cKwbNWENm5tTRr+VkwZstjjKDfmveQQdf3l/Ec75JyQXjZCI4h3MBTL1xI7S6gFQVeOfeMIQCeq7
mE2+DYaLkfs1xWof4uXDgHGCnJXivp6WmTC5MJ1Hcs60J9amzhcuiDt+xNtXPkIpepG/jEIkxvSF
sM8bSI/EqvzTfOy3InIl2Oz8r0GhaDp2ZnMIkcAI6ASHlxF6Xk4yDA5VWi25C881lf/T78QzMJDW
TXZLY5s18FO6qbB0iy7D0NQMH7DWVG5e9raskEZakj3xbdTYtb8alCsZkAilrp7syhBf/EgBZ6cI
2bvAWfX6DZN7kO6dZTvZsmplA0+d/HkY1o1/9JSNHl1GdpJizedMGG0V/+lS3or2gtRUIyxW8WCa
3PYh9KrxLtNPc1OyVuKmok4O6ng/5CM0g9xoWEMzQLo2NSXcz23mbonM/kXSOe16mae/EH8xreU1
tjzDO2gEFqubnqLaOIJ4QYjN7UYeUAUOSOtcoW/TcidpslmYbVCQGlBaLjlA1jfQg+pp2lYf+bJP
5pN9x27YvBwArRganOs+Gc4N1z9aN4j8U6Pgzm5KYvh5BYE0Scg9q/CHmEL2rkmYJh3efoVAHgEh
+nYACXtAV5961fnUhgvAlVpk5JynfdAdBmk+JvOdI594XbpV9FBrU9OYz4jLroAQFE2aOcNCpfYk
V4JMSwMK5+3dH7TzLzGtrVbvP3FPyWdLlKFgYf0+Sxp8j+ATBKxm4dg3+1BLMuWEne4H/bCM0jFG
uIELOPBTsBF8BdSVypTjUEbO1wNCt1MFPo4qukamOR2qgXnfVCc0W2h1p7fSfR5R7KmvRtWy310d
VkezFS3jLtL36WejpNForE2fehTgo2+Z7/d38e2cR+hrlIARGtqY0cYAK22hKTMbCbx8iPwjTLUh
40KZAD+TwzV0M99TO/sE08BAeRIWESADeCudXvO1s5XgdD+M9HDGEliC9u/xTmeMHwVliYAWzVlJ
0SzcJxvrDKLQpCC41eDOfSgghTPqOZtbPDGZAU1Cd0K/Q6CRvBJy6TTYWcNCUS95L7hJWexG1/0a
HdCbRuKyxdgOQCu9YM5J2VrgdzqiNtqfr5TWu0osP0/cfY2GAVP5BgcWiPmvv+LHf+yZNOgPwaQN
0OAvmpTmf5NaAfHtK+ZaqhmmBNTt6hxv1fnI+gPM5wbCTCl1SDUYjPsqrN3qEGQheHm8cFFuOPrf
+gW5H9NKwnzJ6hiWZmRIhEq4jqEKwWX/hQQ9Hjs1mevOHegt79zA9AgglonrERWMKT2mDNyeXzsq
D++CYGfqy0E0/qqjqTiv4aRTfZJCt3BC/dGtTcxx5PQX9x40ofWS/dxhmOYMeqs0qC7KLqLrWjZn
3shzg9v2izpbIVmxMGrUVKK32vDaCEQ/h29gTL6ubhi/efMU/3d6T4r3GT4j6/OUORxFXPR9fKCW
CzycjZUMKEKmAdi0ogxIU745Q2LWKrlPokGE6BzBP2vB89NGaXghuSi74zP+Pdd1om13axrYecYR
Yb1rYE0RSp31xwkyXxRFmTGrcNjdTyg60tAIxqsaUCt6byVXhMB3nK2f4boL85QsvobirGHQdjlk
EEG1lOvOEWeRaOmoNsF15NHEIWqYp60m1zMTV7u+adR+NIZbqa796+kgx/HSB1yiSHo+hZ5Gx0db
0bQADOvHMbzC2YwCPh1XRm6gDuv6WAcKfYpDw89blyKGgRRK3s6Ur0AUnxmnlqDT/U3tUIUwH3TN
wOo5qO9zbomf1vjAqAo1GjNGHIIf9Psp/lNvyX8H1oJVwBtnM9Bo86n/ROSOCOsP7F28nxLtl+Fw
sZzOcFOEkMq2TwTCf+cmv7AvTeJ23vCHa0dowahwmIECo4cZiymYvDNW+wBHmGkYH6G2wS7hIysE
e9Llm5en7mPjHrTlUZa3vN6N7FqYw/0j8HrFav1rcfW81yBaI/Ui9uAA/gU4mHdsWEU3VLFY8e7d
TeQ9TDWx+qnkIACIoorysU2x9YXQuJiPJThv0Y0aDndcX7XGuB3eJV9KZF9IxxTIZCSLQ1tU6d/D
FqZCGw9mZJWBLd16qQsDtvXvzXqpfIw5zSJ0IC1wKwJkL1t9heAMzCMyKDTpRAmXpKiXuMEcf7oJ
2Nhpqogi5mcbJGLuIro6dzrTZseikQWo/4iXemNN/6DCWE4C5jS82cVl7r++pZYtk+5J7TK8GTQ5
7iokgSRNBF1np6v+38qjbZIWGjtRy33iNt8d0b0MeyRpQxARwZBv02Ga9mQ5CTA4t6pZ8WYXDtOu
H6jp9tgjDnCbCwg6n7u868Mn+UqBq2Ppix6moFp0qxx4eVWjNrw7yzseOzO/i2tfxeBBtpEudpsu
eiO2Cisg+LmzCl9orkbsUhzpXgJaTlOzBkI/yEqTeFzqmWjpJKJ8pFPXnvz9C+9XZ7P8BdIVa9pb
MGIWCt2q5v1dk/dwJL3PCcnPGy323RZKIdLclF7p/8F3BWD3nYGTLfajbMo/kObKSuiK1EqdqllV
4XVERcblySuwk0O0A7VQE8WAWFgd8laGK3LdfN0Q5esMmT5Jq3ESoc0jtUyjgo6WIeiGN1I3dn7d
r/056kallNW9WtqM0VzjpFgw6tCX29yY6mdttTAMVlibtH3Ydtx+m3xJleMJDbTIMGrEcmoIt5b5
Rl8kqF9/lOi9EaQFixLzOL/VXJ4KJVS7d2z9bHsbAkCYOQUWx2YuGPN49ZVCbbFpWfJcfDjgbQ0W
tFHz4AfrP2+F5hj7dV1fx5Zw+Y/7Pg9JbYLvctYTRHmn540wA4BZcNYSCCBSEjOKEXJ8fPzW1oQr
t2EM9qy83I/U08Tnc8ATXMxLhf3hOk5iaL3F3lw33AqIPKpgarNGK9Pr3uWGlKmo37/0mYyKsUcp
GZ6MtnNzVqpA69knTINgwh6/0UE6FqQEtYJHGVz0UGhwvzXGQe2gVFJBM0sbd0zs6Ohqe5GLH3nW
mrbULKsJhTDCdlLLHEmDj18HoxcAL74d2Z4jnXeqaNpAiqxdsb1JpCykexo50pH3XbhfUmp1MLeq
oDSM4eIt5MFqZNTtFh/yE7m10893NohcJ7JBHO1JcOBlxZkRNK2ofkxvtU1U/EfFYg5BG+pCkxk7
gl/+12xjLBGK87CiRmaCVksO0XOUkjYoR11LYMhbWQhYJtocjCuQFkddPTkWfe/lhkt5iSdYujTf
Yvj4ywHY+cAUpW3N6QRxLRFPnTmiM2nCDNMMw5LELrLeMgWc0gsMBGql5s+Ez4WKHyrGrs2QvsI/
zQ1/abt4uCicxGRawCiOdnkWLfdmXJv+eQPG7VPED679E5WuLdEKSqm673PgT/UQP5wRu3JlSDCf
TK/lhjHcElScf96YvQXTl8AuhXT891bz5mAyKFOaLm2ByLvuy/OS46bWp/kAfaC+ShOM0JxTYiF/
wUCKTqOp5lyjEjo3sCLu5CuSvyTEPd74bcUTfjnIL20zh68qTzPY7vDstQlPDvlW94MQendcaQm+
evTxbe9LCAbgm6U99gQ6n+coyA0XyY58mmN8/BJNKEDvtoNDt68grdxcjCQFCnGPbA0xBv6CmZUa
qAk/c+wZqf8srTywromep8sE2BLRMCfqVe76Q3TmFz3pbAlRfPWJ648jgRC/Kyb1yi4Ieu+kgkCQ
Kmz89isHEf4wqGLva9YVMZ5UvBOE5y+mf6ImGGu+iU+mRbB7aMEwaXa9PnN5BlaIojj3NBzBmPsB
PlfX7KhfcVJ27uPZYVoAqqt9DlnYnl31xLs5ZtxUZuSYVXfnrMmFC1k0Aq6WeOIfYsKv3egtbfEX
m/i3imIawnJJikPqrRVws0KsssZrpvbH/Bn24txbP9/WztPCQQ1b9UpW23JYh5XaKQq6W2FUos5O
1f0D3XC1hYFBTUd474R7HkupJOVZA9c473/OGp08Fk/hRu6UPjgJ0aSuHeTwVR7mbpN+CJTYpAf3
qubc41Kuw+nkNF5H9vsp9/j58MOENY18x1iFC0mNAlw69R8WVJB6KQQSk8AGRD4C86TajDvoqorV
tO6YjMULxQ4Zf3/9GYzSTB4EGLs+ogKe/r435+5835DUfGOYpfuULWIFCjcNY+3/oHDMy41zlNJ0
SkG6JeJTt7ICUtyOuqd86RHXBIue0RI5afXvPJiBRO1vJo8XZM+SyopE3XRBNZL/tG2cl2EiGZkc
ZLH3F7zLhQzaBVrZZjBgq6kMx/WALz/s3pKmKPO1iLFMpMdL/piAaFszHKvQ8/ql9khd4XNaxM3W
kg6UalA9Jdg0sUYzzyM/miUJKsYc0refpfzE8gYsLXHD5K61lDmK/EGxn1enxuFDXu0BoQK7M+hW
jN4DmlMPHR9FpYo0pagIiyDEeur3kRkukOZD4nOayohwgI4RdHnSZL5BrEJMAcWl0kGxCx8LBA1K
r9NUgDuCELq4s5pgE8UZHR0qkhRL1wT3gc8rI66bCdZQGUFdCOUmklW7isl2cc9o3P7psPQRNuoS
jytcs6ILG6czHIie693ldEa7Tz3ZS4lfj4JKLvffgYkik8NTIhkFnbr06JsqrCXb7c6xA+siFu05
+0SRHSeUWR1iw4bDSUvAyZWdVqbJj+BBYHuTl9n07ka8S53Q7CvIxDJOqII2vqq2S25ZWaZdaA5m
5XqT2m7G8Zo+Be7RdHsL9L/VAEU4iwMm6XJAEoPoCK7D6W2sDsk9zcwXbBoGyQiVMknVWRg5ZEUB
MyNuFJln3ZJutgcYFhoP1u5rIalRzwAB+EPa1JGE1inwaIrkf8P0aF3jzcXegJj+QuU10yyyugZ7
FUnfrmTSNzQ9zP09S7v/MfE+KBO90apf42aPNSl+ZS2BVJSnhdDTJcrZSYN0+yG4lSXEfGNJoz1M
GUTsRUdxkxEHxwNy1pP/wb/39T28X0Mi9+l/vvmZ40MfF/LjggosH3lw938bGQoZhEcx8jkEbQ3o
wYMu+00eO8UJJuppshse3z6zhYnURJtZMGG7PuthUfaC1I82CdeXxlGJpY/gPgcc6JVXWO3gPKjZ
1lLVY7EyeghY0hdHyZYWkzWjdk5lpCPjQrrmQInElt+Lh0sn5Czz/qcpQrUNgE2HeN/eqSoVg7TQ
EKjrN3YA7aoXqJxuv+zwZKJAai7Z22lzlNVk7+sooenXPDNikvP7DvP2aPhg4maQRWVsT9wuwMNx
lvScCNDMI+PZOe/FF4YEE8LhiGY+/M26S+uwgsKJA8nrupRlwqa5L65pibvEWM1ce+5M9UZ/t9fO
qSSCNaGnOllIVkb1SNFvlRUhj+gpwP3g6Dp3eh1UrX2poZk86iuEhJiCXdXwjmy9S0S/uvSaVgeq
J44t512O1BwsWpil+IH6XCpR4RgbpStHSX9MGbud0qJn/m458Y4td9lATAwa5SMsuNeAVTh037Pq
cxI3cFujE+ZPKsZzl0NCVxRPoHdcYWvYLlMU7TW2alWuzjkiuAzsFv6UiO804j7A4tHE/n5b9MxY
NmuSCpAA0evdCSd3Pc9gCTHywRYnsGzYBt0VWRGSBSX7BO3lIaSESSNGTc8xWiCAB2nmjDU3E8wS
AfpWJrqZQ+vZwU7y/rbAllV9RgxPP8Z1IF3F1FKhSaW2fUzXRV3e0pngmZ8HXjv1uFnrB+nsuboH
Z2dyoYLr2JvqbKABzYUW19TpE+y7uxcsWkzUU0FPpsAN4hxh8lg+NcCqGAndZUoKsV3ZzeL5+Vy6
I8p+a/0IVSJ8FZceIg2vekuHWGLu/meFoA+srkDVT6JW8O3DUuHdeeLkqwrNXBod/I4Y2x2Ekkg8
Jv2xTQ102jlbpxq6v1LPgrkc4z1x9peAbbcYR1oaKu0ifYVmM3oDxGP73Q+j+6GYjy+EFGuXdwuA
xc4mtnoCw8Hgf2GERBGpBp9KcLT37jlZi7K5JPy+idme9PRWa1TZzifByOdQR5Qqqn6utgdh3dWg
yF4DGpw7ucQrD69QKMfaPMl9VwrWmgREtqqyfMZhk+UDMgBiNapj1acNcjEKCkZ9B/J2ZZ/is4Mv
0CmgwSm0e+Wr1yg7hVFdy5xBynuGr86ole6Hjhh9YLFAfzNyZTmlU/XO3D6m1/Gn33E9mLyvaz0H
ihUEkwZ4aWu5EAJePPt2KAswWdcecCaXcK/nZoJpU2oNX8MO+eSKYv+tFL6opUd/6VTKn58HOOpf
Zkz/5N/wGJVFlzst+8iCp+k4fYHmD1is9HGZJEJinE67NYlTdpD9od5VQ9W1rOLmcNn5ROkLO36m
Rb1eJYEs2HI+jAmlzeotGS+Uy6B4cO/YbzS8OtoOtLtTUyk8oEBFPbN6W8zSf8DcK8YpAQe3leGV
2umazA043M/pfhDNViZLVvSeD2JH04czslzomO0kVCX6c3BAWWTL+5oocziecOYEgAlZlfKoXw4s
e4FS8CwOA4qoMM/TIf3FB8gEwHVnM1dD+jntDdpl9TIfjKFsl6aFhsa7oME4yrlQuLrV1n89HvKl
WstSZGqfu4qu7eolc5kUqUXLCKdQsjcuWMdIaVNHvzzX2q89AyCTewHt7PCCzD9Cr+ynE0m9mncC
2Rteddr8e1LKQvBepoZpfBCawQnAIxiszL0E/X1mGr6hoLgmrX7lQ8pr71AIxE8nVV9oiFVWoQBm
56/WjJB+y2+OdEObZZgT6c3iaK/cFhOaOOeR74HhSeij3FnraR/dPcvFpkcAXeLDAFZmA/IbwV+f
cmJHdQBIOJCd6ui5bgFCXiAibZT+DO1jpGfEHFWTbOTAOAIWQc+2PIeiCGq8jyGL89o7P+OITnTc
uGmjmwgNoolk6cr18kBLkFs5DUbW3+1taJnPH9lZWMsbV2fJP0snTZbYU8CcJfZvmzmqj/O1J/QQ
fkbdK5U8pWXCVD1HIP7eVOW60wiHSi2/xRAs279vo0iH95KSurgPP1r0Lx7NmDbch6NJkeO9E6FD
nI/flWpC2lQrphrp/YQsY/zwUwMDnTYq0WryPKDPX7wyuwy4pWrXC5TyJ0b66FE+AIeXhynbS7Ti
w0vhdgRcG6emsth6mqRjmfG+95p77nj8EO5Ef3x8aKcZOL2HpfqTpWc0H2opnfaiF50LqxUGLOJE
jD1S+DDReL5QKm2GqXUsQRiPp6KXC5bErqEaTjT61P9NICHYTtry/POqbhMQD+MYd+Vm/XZNkIMb
Y+2m30hbmelLc5vj74xvuVsQCIr0O5EwlrIOyS6JD1gDrCA9N3AgoK7HxpUbCnJ/CmWSg7qfdRr6
RQB9rp3GKhCpQkcg4OqEPDrqyzV2nItC0RTMY1KGflXMl0tXgtA5ZwRcnQmT2IOXCSEmleGqkRbh
e2OvvtEbHqqXlp7CctGg5o1jzUFlUf2XDpn9xqhswJoxE6wGYOUrP9UBvaPctgPVlxu81xzfFXoM
8IJb7d76Ni500lUSoS78DykldM5QvNAhIPJvCbtcY5E2ELDPWYuijLcsxsx551OzO5XUsa+1AEC4
DReH8EdG87h54/2XW3cT6mGiJu6dL0HUNiWR5PqWisHNrXIVCPd7WOiq9pcDLdoktynAl3hQ9E+q
48WjHAj+F6A/ET4za7zE8mA6M54/lGCFrplY6O/m/rPoZpW2GtFgHo2C51FZc1lxYuMD/jX4Nid8
k5SITnE5yKgngVl08cwjlLIpPgNZ4dzmRBkOka1IeN3YjvI7Hg/+qJYpgXY5JVuigDH4b9YAJ8oh
PGAcixUiig1cnVfLtK5EhoHJT+oAunmBSQJFqrShIFd2BP4zNxQbWT+wNggrIdd8Bam+PVfZuDya
iEiZcF8+kNbezYEriNr8B2Zm10mCyYJUpqRAZsYi61VYkomWRkRkZWPN/Wpy1aLaOO7ckrLigpXT
al4ae762tJJj1Bn3GV3jVODXvEIa9H6gjqQXddHFl0nTqq+U72eoBaSjg1rSDdJIWp1+PtXJDlRR
HaZDEi+0GuQgIDH5DA0VhJwBlVL1q3sb5NQ2ee2mh5iUDZaalcw+ibvl/4+m6g3qfXrsqPZCvu34
fvrm+N4hSDn9DsdSzvabYPkyrAwzCohguadqVSk/WbnEVyHc5IFau3JgpzRa+DxeQa+ckOzE81Dm
QRlaFURwpNhe/PhIlycpa5z1EWAxXTSd3GKq4Uw669obCnQyUc+WRqS9SBc80GYFat0OLDlW9fOr
dop4yDnq7GZ3e/PLbCUwP6lx5hDAdnfJCjXZHh7DjsfWtHQ+bvwQmAPDz2kXRMzMrMbLTestsk+p
KYX5WulgKrMvNV37fdK4JrA3EGIyNiV4Pem94mVkYpZLCl/vV2JdNTUSoErDXVydQ3BMR6aW212j
/4y7NEyHikDkNKHD93Sjs6Z/217gvd+ECAKk56fxpbwkzBzLZDisanenqj/DFD02f5nw/ikKVeon
6z5jvWg5DDdHF4yoqcFt8yurENxpkPszsq82CndeZamfHzBg/d9vsFsknD6284Ro+ljrWbguOqMs
GOoQAiGQQzz7j8546Hgt+qII80RUXAVA3bEiG1RD9/Iya+iN6KUs8YNklBDs5FozrxchKmqPeAOB
eOtCY9Gylg5jAvujvbtW/CdX02DVkoe8xZKGbYkj4TovCV2E7MUqFQgIZXhSSdCsdBP67STkdut+
E6j1lXOKZBN7PAf8+vy6gs0ckxk6ia0E9yVuCp06E81xIkiPkyunEJV3rs2Ik92UDpyTEB1VLNrR
jtk8inqlN1o5VuTf3XQCmmxxnIGUYxGYTaBA5D9cwuAp+QvDLrAA/salLwr1Bh/2l1YdwV4hee4U
ThTs8DXkE51MTBbmQpc6Z9snqFDKeZXnQHKd0FFTk3/aL5YSIfq6dVlAEj3DwpvJ8D9cPmb4p/1s
Am7di8wzaE1n2IRtNt8CnomeNlXiuujwVDuMCE8edpcuHqnB5Pd6w2WRykVadG2zsS1WfmhwYD1z
1GfFgPFXRRStCGNgcuKKcjKm8xdwF65lV9N28LYrpfdamaw+y+3RnILoCb0UMfzDuTGShDmWqJD9
e7e9PyXQ27R4b1hPeZw5HeXTsx/AsIlpIrXa+6Pv0GCcXvN4WVrCD9msb5Wm+K4TNCK7WRHMEPIE
PeD+UENT0E7Sl5xD1+ehrQ88wQ2wxDxx48+WPwmHQRp80JnpVfTtRSuD29xTlHJJYU9NgiN5ESQF
Uuq+P1IBRYkRqw9XnUFyHIt86Pr4m8k+ut8kTD12MuHJWKqf6eeCyD37WO3Z1GPd+eZoxpyfB0UC
IpvLbu3G9QhdoFAwgE7KGyFdyhnsiHc8OFmvwAH/UVBUV59TQz+oo9tmuAGDnQNq9rQ7KiLJ2l5k
nniPESY42ignvaRo9knJ7iFu1E6YAws4owHGmq+J8J4pPllcx8n2aBEGPrlPvKOpC63DMtvxQRNi
T1pnjIV10RszbV2Qm0LSyToBnnXRaQzXJU+B19Y2CWmvOm/DzNJveXGBj0RbrPfL01PjYkhoOZgh
bEYNCIDag+rOb3Nify5Wy3CAY9sYRUhRkcdFIAIKAN9cacqY0sEFhya6jn/dzzhA3drwJRgxzpln
1ueqN3Yg6mAwfNUeJgRe2AJ5EFR3vjJelhoSzo1fE07wI9lOLAesBDbAhL48APSkEELY48m8U/ca
SRiG4zCbvsJieCLt9kxt/gLSUXeurHI+a+bMRVRE1RO2peIoVYZx8eFMVfPED6EhWSXUqlV/ZFNw
pRtxUnffZwkm3KG3w9rqu2o6k0cJo4J5UzvLEB+8MfoA9ekohudTGZkTLetGqRJPy924WOhXWazT
fE3tTFD16tk6M5EiXk0C8dzM1BPKfmYKTQ2vMMyJlJ1voo5J2Zfm7GnRaPFqsCjDMdJMoFoMpgyg
M4biss21pHzsSTtcIyf4rchN+k2og9861WU/EgSam2xVEuAxacGcpbmTLy7339DbPYjZ2Kixf8MU
brhqmOT/6B77EvRrSgVmVamZpwT1PB5TaCph5pF2bzx8ryT4mlAEuOcxjg8BlCvMw4ICCh+ar8RS
y+N8Y4AKAOqtdVZDkWNEn+d1iKOPsg+97nG0tMLogG/QsmJFBr9lhBu4KbugJPw27ylHoElMH/Ed
DfHfVGAJUEDORGyEteEKoHCBFDpu6MYOFhMIXoW7xlPLlKRe7Saw6HYxJwIYwptRNL70/sLVjKkE
+oPeKOQhRRrhQioa8r4YVlO9K7AIxv6/+aKYywSSAYCUGZoVnylXYukLz/TKk3obQSJrkHBj6tcc
bh+YgUgWm+a0lHqfohORzZSEquJG7Tdx088gTjNVM0SQCgn1eoLCjN3QOBRsl0HfJoIGtKUlVYrG
feYTTOE6s/LFt6n8XdBZw7f5/hmgFFqYvLXIGjRRZJutMuvoSYmvpovrnik6J3YE0OZRSSr6oTFt
GjuiuEIra3dq0ipHd3VtewMSQVsl/8pDNL4qJR7sIvZdDo6sEa+Nner2h6moHwL8huZvedeULtnw
PODl5g6JyPxIFG4g11JODgZy6V1ONq1dvUsLotE/c11JQ+z9iB/d4CbaSYGVuRxcApcmBh+mCvgp
d5ye9Bhub1ZA3NQgXGZWHFU6HaN/INMF0M9ex9J9HOj3AXQxEOefbzerC5ADzUNuoXbcY2jYCxZ7
mjXu4+ZgQ4HBvsqfXU8ysZ+LtRqSmkMoMInDocRNwgA0TFGXZTOizbjtTO+8Vhnw2Ri2e7zZbd93
l0BA378drppqmFtr02hXO5gu/VftIUeXESA95D4k8vfXsIGuyRUv07hpHfFnLyylxBr9SEWljvTJ
JysaAGJmsLu8cTlNUEuqEJqcZdAiaHR2NWsvG49GqAH962OWJ9l9e9BrYRhFuQjImGZVv94WwB0F
3M9RY6EP1tkql87YSrYMrx6ZpRQpL591lJmFpzix4xKKKJjckq6TDZ8utgaej989D4bGkyXmlpcq
OeIF07MrrWxOLQ3wobBbJrNnXSmpWBUvGwORE2xkjVtRGacoOzCVLV06uTiRRG7ao64DQEleAwan
/EjyD+TjK5GGQljOH5i+/Ff5D1BmhoPf85/X+05joaNswz6WqO2a8xSJa4QKRL5UOec4r9xpsuRt
3U3XFySDjFkCgaT33CNnE/+j6yJn272wMRupszwgjDOB4JwSgoPKEJ+ZTuGY0h+rYSNLJqZ8IZS1
GX+JiY6Ultl1GJZgzUsf9CS+iHsXNKbesM/JC3njtvK850HK/k8b4OF0ceyJZx/v0VyJWVqASb+4
l81kdfFCB+rk8459V8OS4rLGLtor0C/mYnxHYqCarBsn0dNhUfC6dZZFC7Mdgg6KAEYxbj10G8FR
0sxKcrXYUNWeBK0Hp2cMiCLHXkQWl0TYvk7wJ0rDt96Vbixd8ak66hfn4uJbZuUnfOwxshSewxf5
0sYoaEIW9lwkBU1kJjiQ0FAc8XBdrrFZlbvIknJuVgAafhs87l8MyNJzsz2oGUD9Sk7PR2zFIeF2
XQKaYD5YQBNdusbvNZme3G050hU/IYbY34WW1LDLAGoO6S6yallgwW7S8tj7dY3ggT/TYfbCx1AB
hXEGcZ2yxfu76EYAm8dquvmfj+CF0CpIw8AHDiPolV9GQCMmHCSsY80oF0sO9Hsg4mdmbdaPDRrX
NEDHS4OkEtauVwcs/QeDZ2RBmeOLDHmp/5RqadkIC4OHixyXAs3ih14DC63D1dPyqqJ8d6kO7DuL
5pAOuxRrszu3ubsmGOvlH9wpoUFUecU3otHEGXgXNgC9Ci84l5gBj87Aj+TEOwBFNssy/wD9kmVH
tHJdkCp/3N8WRbq1/P0jPLbQ6oADMVulkl4JCIZZVwURMrvo/Gufmyi+SENfeYFevyoDqyH+BT52
OIZu/F2+mohyGSwOT3SU1O/4ylyrmKAM85ZQ/5mGI/dld24FV1/JmW2EHNZSKPq/lU2CucGAVzDP
mtoR1ubDhl75M3ESyIUlQHF/zY5Zw25iwK4rqqmzHlofCyBG3p+1WLei2HYVUGl+R5wXnpIw+luL
HGFUbS4FIIC18vIJQ73G6BgB2WEOkbT/zWL77uZeVwYuYbAAJ9DxW0E6GdBRj3rLdgGqlOdguIlU
s8uOV8AI+tToq1fMVs9OLM0BZZKE1oITNhDru5ejyGrVcj2P1LYZx7ice3c3M3ayr4TEdoilGw0O
rx3upx/jX9XvAD+0TXbv591rcbf7ydfOO9vI6T8QSv258QC8THLPmV+nw65CElidydfnv29y/IRn
SH9FYh1MI8C2bR6zIe4B+p7V8h0qZmrb7nIVBxLYSkTiMuMlq1IWARyYtwy4pVXkrkf2T80IMcNw
KMmdyBiJZ8y/VvqpL2tmobWsDe3vFLg5v0OLYaSbFTte+eehcHaXEFj36Vi65bgm/8KFCxcjh2nx
oYZZQmDGjE6qBtkdKrPZ0dasCFPHqM9wP8KYdZR6lGH9w2Zmjj6bi1Fi2z7nxg4mi/N/6NjiZKXz
QFQ9OYmONzdQBPLjMQ3rMQqjdw0/zxOg5Xt67HNFu7WdSTrOzO8ba25jTayMGJEQTkrmTKXwTbAD
edg+VVMF0jylqgkceGQCitkHL8tMOs609DH9ySsH8Z7SGbssCluC+DXXki1RKAiFoRN5a6Rr1y7t
JsWXMmGoAuirsMrirHQx6cgbaeQRVdRn6uqBbgVFtNa/cJJ6vHx5exCDH77v43In8Soqlk0/3bxX
rixoClxieosIq3jTo5cwnmLfajqh6pogq/vVA9fzO+cW2Y+8w4lLqQx2ahENRIAnaLOwNV40rByD
/UlCnlfapSctZk7DGIv65DIZoo0z/xb0l57drdMjB3cetv5FVUlubF+gHodVlBUtxiG6gCy9J1Gq
43N/PkppjojsgSU7LkfySUlpsdZdjt0t+fev6nvPSl3NrJsriMxIV9IUFZpIwQvL6iy4rBE3mZsD
HDCnDO0+6xPdjRYEB70knyJYCrXL6TKjkPjzffqHq+mukTxqY/isZ4DXbcMI4edWQ1V6S0YAWga1
dq58MUi9oYh60UZy5rEnb8Ysg7h8Er51RIgXr83iCEwOEXQ2fLJM4Mxx3Cam2LHoGLcXERnOGjPI
sU/S1vTsWdY5iqg+lYYJvjfHX6DD1aO/QhdLKcVEmIK84zaWQ9LaUOLfzX2+w3sT15CB2eOdTUTo
ZH5i5Z8/mrR5jgRa72eDG571IxfnrtjQnl++Ex3UmlgJ6NfvCyj1AoqtMG8UJN6o30/Q7lK/Zo12
RZBj+PB6oWtWey5xBUDW0NjqM0JcJFCgm4BMR+D3NAfP9KSdcY2p/xikqIhHMm0Rzs2xGFspet75
MLFSAqr14QzPtnLoyP2SNLS4A50YH1estN1dTeDuN3reDapMRToLxTG9u7Xw9WiZNhUbIkzE9nLe
td87pPsAY1PXOONyhXxiqGgBN4x4iLoj+9C800yBMz/ht1SqPeMhLTwlUf8+vJn4sVJZNcaT8qVY
5HnHVLLQhw04sI82Lf9j9dp9mDjwJ4FRlWotXJ1OqiqXEThXOf+6snMS97Z1A4oMi8uwx2Io2sUv
OF0EhwxlG21kQoWQpdmD2LGOspfy4Hq+8szd+kOnQqVsa3nQz7WdhhxskhnXEjH8UPLy4ScxUM/n
FOKYOQEcF++dVq9paoH18EFgtyf/rLGWGMmuXKtAnlzutPmqzOOvi0nKAWnL0nApxUOBxtT8OnpM
9BscuQWDtZm6blYM+9RJA6Ld5K/NeP6NaS3ZJow7Ov6FQBZI7wuLz8IpIU26zm7kEi2HEsTo8cyJ
o3OyQiTEn6RFD9Tlntv57h0585o+E4W9P7HKTqKooOmq9Nnr9heZ07mpWJ+4ssM0n1TB4n4Jq9Pr
HTcxGEOILmuTdtjiY3T9FvOJCF+gssDLKCt1R3wLXtsy6Ipw1Y2yiFG8gBgZuAwqi2wjORuz4EYZ
OBOCKMoUcgZd4+PB8h7xrnlhMkwfiGvp4/6KnfNQErHnQ2KytVu73okISLIYyZlnTX4fROEoOLpY
sGWrrE6vIAaIAbA4T4VOE0v6UVp4i/uHTPeOA9E4yJAT0HxaMTSOT+TkQlmQjIvO8wB3ikZwrPQp
1H88LGN/Y8RVi5naukbfxH+k9ZEikuJTbtUAIubxwBSHHFimp9vOgiBkgCuMXgi8dLkafNwI0ima
8ZtOyrS7jh8rrYb2yqY5q3L/xnNYroUX+3FMVVpUJZPjHZL1s9P9gDV9AzdJICApAtJxCCNuRF4x
3D9lYShPcw4U2nuJ3Kv8gR9lJubsi4lTNqfdfVNhGKeQMEAVQ4oyKQ0mSwUgq3mt5H8lMNgvKoH4
GtaiZ1fZ/WhAbYwNclAqSGk8AtPdEvmzeNDtbFHwUUUqMGWA5DFEJFrvi0vC3dPTbo8cObgxXJ5W
GTPMIJuUtDs0+2N81bV7DJCl26Er+D+e89wMfexyOtur5uWyzdOfcTC1jKs/+zoYBV4mF4XUdV6S
kySJeWup9n+BvBTeQTBAa28g6MUt/PVi83JW+PruK6aLqpMQMV6PbM37nrxwx7eIsww0yZT1krRL
o+V3DkCzNxfZDfnC3a644X/PnmNjPnvDQPei10EKWGL3/jB5+hfdsYZe76r42+1uPFUhdFkpA0N4
o0pEtq52NZ3cPXjOrV+MP8MErbbBIKc4Gu7iqKyEMaLKnT/R694EVYPJksITXsdKg9h8bQekn+C7
ukkEDe4mU7KfXOpG2cQ4X00XNBTOyAoVU+TlgygrJUqIQmal+b5S0RYRy6BoQYHNA/Qc6tu0YhTd
akSTy/xWt46FOpzPkzEDptT6PMQdLKBBydlrjEa17cXzKlllx2OSIoSiRvnfuuCRSfi1KMuntrd2
CxP5dA4C22hR381wzGaCgPyd/0xTWs1qgOEWn+2xVnU8LGM3xerhDfYiXf+MBppN8GRB5Q+AQzRW
DySdDBeR0Wth+YgMjTZ37HHJbb7ZZH7VWZ6hz26Ufpkvq6MB1YzR3FGsNi5izTahWxFfyZTdv085
dAYkUhuig9qYfxve0wW/Fs8AMgLIX9L1aIHkzk652Ut7t8Wtz9ELMVOOcAmISyJcMK8badwJyKhd
x+r7X1WtwaqzGfAVYo72LA77XmUI27MGhDfPUc+GTA1CZ0o6U0KFrKob6GsMvA+o+HMwpkRRbywV
jJPzt0x2ENO46EQWVQVHdloEJH7yupaYzV+im/kGfUzu5wiJEMCQ56sEXBVZf4CdwcGSAXBHxrWx
7RG1U8pZSm8wGUsvr6hgDY78i0tVDvpQUKCdOYBZk3I2REn0N28ghLZh0dwZQkO15YOxam4qkN0q
5cSvIqmxlBr3gHRz7PaAdVpzxOFbM+ol9CX8jtwCcUHsX+znbpvGtLmITA0Q2xB77SSA5DdaWgZS
gGEr87Ve3JURv1gQULD/LgPvjbRFBTzjoSBJKjuOodbYDdNwGzEB+lbetJEHYX8rhXhUh28e1s9k
PG+9W4NCXY2Qt7Rb/yRgJtrd0DbE0rVd2MGpmcnHV3/Ea1MCYn6b51XYEBrrTOJ6ro09YrRPCvPh
lAwFfHpz0ue2QHhu+TI4fyfuCIJ3WAXs+9oGKXfZy0R8qXfoAQf0akEKbpiVjtuOZEHYck6PrT4l
XhPqpcj9tkF3iw05K2Y2K2VcmibFWx3+hyOg/p3wFPCxd166Zv/Qu8BQuODuKh3MXh+XCqXDqGL8
/ZDr8FzmfkVMOk1MRYyytw6tu4RcAAqJOm3Dj3wKoMDSB5KW9U+25mqeQIaUbLPYJN++oLOP8VR9
vh/cnd9zlfo8W899wGEtBou2rVxMsgu0m0N5OZtiLzpin5Jp0fvZ/kVn5WWB6j3sD74lXNj3MinD
3F0VMwl3RO8mqhsfN42hXlNRA3LC/IM1iTDGRVlsab809+oVjUeE+iI93KmA840tiTPsynkOQ1IK
B89XCZn2PQ50Hftc8kI2EsE81zCuqYkujACYbqPC26rohINNrOqnfFnvCS9lZ4n5BixggIEKEXF/
vdkp9EEo+krjT5LtIMCp1zgVKmXHbePM/Vo+8uAECdJMzjLOxX45SA2SQaG9aKp7WYFcmEEq0fEw
7lB7lj8jg34eTLuEPe2exbrx9hg8D3MOCeozCtZ26KZyWJQfH1TynmK8NM9fPIGL9Lvghc31dE8n
VleSXZGG1NZnD3O06cU48F3GQhLIU3W7XPssgyhUmJdTWC1hzzabXxs6t8Ywc6B5nvioTHHW5pLI
I2tdZ4vaueQmcJFrIJkeBjPbF2YfmmDfWwpn5fT2wBPi4CDU8y+7NJxUazpJj0I9Hot0qfF3bsNE
SV1T2BPMqQb1Q4TJ9FlYOrH08oXhaey3IaoZtfzbONB1K1uU7ssM28BYySIBRYqrzvQF9cfKVCPp
DJY2lSjQ3JypT6zOIsdQXQWWSJo5tG14vKb44P0GevNU5gbBjUcumxU3CA/8PGe5bLFcRcuNt0vk
pPQ/MRAf3CXHaubxZfMzJNvaI3ih4zgx0L3/695tdp8GgDuKH6j5piKvEqt0N2ALFEegOf6c5xFL
SqiXQPWQ8GSEybS23fJcKNfdwOy9C3QAbY1IjHXisGFhk5IUtS0ARNoJkymiK8ZMAjYg5LgpBEjB
f10ZWw7AIVXoUPHQrxZW5YqvGPRQTX/tRMUyvXtmDX5+0ptoeYGWjNxvLa8rF+4VGxYhBGABQWuB
080F2w3tLc1eXExWNr8+ZskTUcf3eidSvb8fUfPSV/0oRdhc/2xfjGDgAoVUdiD2tz8ptZhgACC6
+LG7ftQBqDfjUXJVy0v9VwiLcz1fH7EpzyQeUKtXIAuilzbQ3EnA/zb0h5BElZk8wAk472r9ugmj
KTWQ8AiPOELyN0CNssa5ATLtCG8oBpTBlQPymcxb8L7tyuOilSfSfAySO+PKgHq0UKOGd32lZIWv
KsyOEtY736x0lEoT0BKwC+nBPcx0bGeQE+T8Q/4aYZIvSoCCv+9ukbxbP+TiCzNNwTPAnalgGyxg
w7hvQ0b+jHkvWoMwzpvD5nqhDWXw2H/15sApj/ixEX9pK1yD191mITNbhVRX1HygjeECtoDyYWhG
maat3BM2//1RDAPem+EgAIwv5psSqzQOqr/huHqdExBRfJLc5fKkKKXJWPr9ZORVUHl/LFiyhCYs
hff0f1DfW6SipDfA4LmTPGjhPqugikYYdOgJgufZNMa0zZYF/A3OZgrdqwBAEtQUbT1D0k+r9Z2P
5pXB/hOAl6Mvujkd5wscqY+9dl1m3Hem1ddn8X9at3h3ktK5lhsp3Wp9yzcWxdyWo6bMQx2mo2+2
XbRvBt9Z8V3GeIaFgoejV/VZmYV50WJ84W/Wb78LHitf/m7EEp6FbR26TAaqwcZTTJbxAJpo/oam
xofPEu8+3UAS1kYWQhr7kNOrEbIHRcYx8DTIXKkDDc9f2qEST8DOM1zaoRyrte+zJbWrjXdGrl/f
jMZkqhzNmQySvj5qI1j7GxvH/iwPT8kzVal7BbinmAuSjMV2Z4vP8O8PzIEyMXQ7evZfT3Eov44d
WcEc3VDjRIHQJUzlHB5tV+zB4rp1ZDfGRFmN7PczYIdpO03M+UACvWhyZ/zvHnBXfQG+vTOnvcVp
VZdJc3fRD0ystu4lW6/m/fM+JpkQMIZnS4jwZfV3zdVOPqCRqhp8qVCN3GQsFiyuixJRyJi4vN0D
TXaUMQbpF8mVUH4kiaFEh2kzJii8meoe2xzuDSfUD/7MpwubfVynhuRx3YrdKjJjfMPtk0clwiZK
wDFsuCW9/XqvN9gjmB2D82GyKOZBSXMBRjdod/BGNI1fdnWovXrjJT2F6e/oEp10z7CdKhjyyP+X
Ny/z4UShq3qE0zIf3IomBj0PWNGFtwETessDbFJ9hEbwTjSB998gnX44jHR17F1xeRzpA914MRqb
HwSO3qZD1PfPI9Nva+K2G5rt3WtC0KswipSsqf9cf68+mdI/IL+Ecdy88pjaRp9ky88ElDFExds4
8WizaM+b6W/1XQ6AmTPYnpVIpsi9wugFUf19aFSDZsfMDf18jjpPs183K8UPjhkBFXbbSFz6kgL4
TZ2hwL2+l8geksug20b/InuYRXkAsKC//6Mz+Pj9uuCRVsKSfLUIeLOKEySPvePns0D31YvZ1GjY
L8HnZgL8oRLIjioE2rJneYRAMpbYf24OP6+sFmyCpiss4Ad0tuvaUqLcPVrvVky4f5wKDi6aNfPv
Q1liIrsfKk6qwQ8eCZx5mUk0ZVeRWZKeRRui/8t0+MYYdqSpgcBjxaX3znk71aTBwVpe9vAI2/zl
dy7Zb81o10CiVQrj7FQmpfvRrUg0WibjU/IUdKw6nClOh3gnm2RvSP7ovH7FP6vyTr4sWYijhcAH
vF6lxyU5ZEDqAkIfnmWes8NKcrObyDgN8dHnL3f+mFr3S5sOhHVWf3Y+rB5tQMoOWufGXOjtser1
FFFQlQ2CwhUUsr+xWzrHGJYKwNDzmEazU6BZEhJbFK8x5L8U72qfqkhiIZXLWSCxZ0eGQOTg+A+s
ZR+sTVMapD2eahKeUzXqgfBNCcGEN4EeUuvhHuOC/bP1lNG1d6XgJdTzLy9cIThAq/iM7Zdh+QRf
dn1wREts4f/+AHTBHWsAip8QXBiwlzomEwgaq3poP7pH/q2GtZ6jLFq8QprM844jEfgBXaRg8YsK
EwM4LetFJbm7AV/hP0B6g4OIAcuT1UkGHIu8HV/CuZtasV7uVy9s96szZPJGfiuDkkvoL8lt6DCF
chnt5jOLzV2RsGexKCt1i8GttANcK+NOcMPdvg/Bqn7lBv/J5uNN3COPlhnh9ra9Hj/WWL5rW9LV
AcWVb+CwgyKdaMKdGsdkIuWQ+WLjRoh10Iw9v956+0rjGVZONKdxreUnKGNzsm7dU3QrUnB55vVx
rAcZXD7r0kq+BsMW+Kp6W4fPa4LK2K5Y8H1YAFnDXkAfxWK6IRzgef/+WPKvJ5QDhl5bCS5WB3Wu
mpGT3tIL2HTNkOyNgWizqQTvuQXfUt8wObORLvlaYGy0XDq7lOY4RZumF0k9ra0bHqxvScjE0lNf
VW3CNPzFYnIwV5pWnj+kixvOQc8y1Vc1pelSTKOF54FkT9HJhbrp2TvjD4q4XA0xgh/Kbdu/qdDu
XDzAJnDtcGZdXTwEniRWV2dwHOdiIX8+zifHB9J122oFj3Dfzbi2lG7QuxRO2iMkBLXxj4gU6yfM
Yo00eWFn3Wz43sAgpTHmqgyCMbrxmqIPgp10ePkDQyS5FuIdCvRbF7ds+ms3CQwtXARbOjlhEuTJ
b2/jBBeSLJQ+NLaJeVvcP6kp/R5z2ouuVc28lqG1Tkv8ubljHlZgBLH5oAX2OFcTYcO5h/POW7Xy
Su8mLBUfJ5HNvfOYhDKkiCKxUPnNa/a0jF4fZSqAVWhbQFN6UelVOp31+cEmZZ1n8Wo65y+PuC7s
fSmNL1YonJz0hddZZ21fjNSVsIcZXmmH3pX0iv6eiosiGhDZtklDatrchjyjYD7gkCi+v2tVNGW9
PySY6cqpGnYT4pJAcGwa+iN4fLp+EeDDQo5XT46V9RfqFXI2Cme6yTEYt/b9Q3jv2/i6OIKXw5DK
XF7fw/Dnemu2AqBoL2h0VLKgH195o2wqKY08HZ6kZ5U2SmphyT0cfSaZWcAcc1AMUQEZ8MxJLPRx
Cc80ujwElE+ucoSsv/w15q2f++5fFroSEQKwAM6XUnNGan3z+n9PAU5XcvPaI2nb/knAXdh2h/jb
Muz8pVEu5qX0qLE3pXcm0R4NWhrQqTvZ6zWy9jVoet1KutZFFWBMD2fyQdlP/foPPthgT0O1GuXG
KAZz2LZzJHsibGR0Mpr7DCo0igyEA6D3IWUCHXbdvs6XVGpRtEtmZUF1Giw8i2feIhfovSTXdVF8
D5M15ZvnLtEMgMxDVcKZkBgPbVZf+gmwBJksOeTHgKqdZ4UiZfbDE5xbPl6LV0MU53+H7K7y6xfl
g4wTymoKwn8bwxNnE4r0IDsz3Y8xhhMAoHln/bOnrSMveijgB6N365D9dxkuVZL0FH94ozVZLYz4
Zg94rMjhaLeIn8Hvs0W1J8Xl7/cUbF9Yui2dNdhI+S8UOoYq9UXubIAf0j1XoCjaUPPAbTT3VYUl
ndtjRTeWznA/BVFK8NI0NMQuPZe3riWqRt7Pe59Q8H8UEW2jYuez6JnHnb2mM1r8eBfgNRMLnPVn
HfK0c4H9Dy9d7iiLFF5DyIvFBFzkPovtrsm2LUh7byCjOaNVO7Nd4TXQv7Usb8Zm37tQqxEb4x2K
qx8fhlXi31AyYHi0YX046Gn5DyzgofABoo33lYu+Fyqqox+d3k8BOqAql5gDTS6Qssn/a+r8Z0zh
9bbjFKm2o76rFN3K8LxqVJsWWbFiJJoEJGFaNVw3VDcc/PK+drvl1Qb5w+n3RTcQ1jllfR5SV5Bg
ohkkWgN1z8CjjsS5NL6BLerWHx1OeceQTLES1L+/XohnIdlpPcQGjuSpZSEyli5+NhdxJszlpX9s
RvWMj/xSofT3gJ2Cb+NDS0KZlAXSynLmb/YoncjqkDy0X7QyVt5XoHX7V7kGKsp6y+zca3Dd2ifd
MFJYRFIUoR/JZT1hOQ34zYl6nPCShWtGu2WbZFmQEh+0+bbng5y7lac6TjbTE+dmOyKl+w5JNq5h
CBZmp6PurKPsfO4971hY6m9cqXmmT9gaJDtb5z1zKJjGL2O8SMh4WwtN52JsbzxSddJBxhc1czAU
B4i7bjo9SAhC92wqInLJl8vxH2xIaZLEISBT8kS2UrcVHtXZPx1s6RERaAPmlTFJyGhMA4tIYfvm
uQVTnZxKJTkAU7+QSRQS32zG521EXfoKAxxxKOJCRI52AR03EbtIvBDElPGod7fpoyDXkl8CUw9Y
hSjIHZ06mphoBxUwQB/GmOChssKdICEgSC05O3qoYhs54wviitSPlsp2S1G5P0cT0gMO+NbWgc15
wP55uONd+Kh3isySAOafTm7HBcXgUbVUyZhWLd46quPpdnpgw44u7BfCtpjiE85ZU1kOkCLCuOxq
SSzunmt/NwOixgY2syRQXABWjr4qYS4IVkceB+8G/JyIaBCvsdeHUiqIlhYXq2WHADanorGXutlm
ElMntqCWg5CPAXQRKs6IHhkNL3r97UTjPpx7jcIzskAXcN+JrIPEBSZl2zPMpc84dlWqiwBwNczb
hSzL29MSvjG0LqoyeJqwQsh8h6I1lQRVwPVwdY1CkBM7BG58hOfFHMHMUyVFRgc3xBdFVtnrWhBT
BvGMTZInWad7stkRxRjLQHvV8gwzBM15e0/4gSyJ7oPcgFscPiBq8jW6Fc/d3HqTzSc2WBp8YB6y
e1fUwEAG7TlWkB/gg7z14wZBAn7sU5m3kd08ZF7xWy086XKyqwvWz0ewjOkoKOBLlrt8z6aX5mjc
PMildJ6WhmrrGUSFccFtc7Zhrc6o72hOpKrYveISxj5WGsQ2Y0AUTor99WxqbJN70j7GcVitBXdi
erxblhFqgleWlOtNBYoFemKID3+s7cEoczlR4QTmJd9Wq85/EWqg9mG+G6Ry758G43jUl+2LABF0
ewc3WAQ25kXulTFMjdbCNfllGLXymk73FPQ0taMmXDoKjHBxXM2mc3ou0xYOvoNwH+keiAs4lecN
W1NGAk1GZNjc04hyDVqHUKDNLPoJE9c/16ZOEsRJrWTcSdpZ1f+l2UsKpai+D4LZlD4UjZ80BlU5
r3BImWL7g/1DTUtnO3nevduTgdizYjBN89XvdgFdpXBAp3+2jrjKTLByoY7r4JPUvp+lic5ns7BX
xlvlBj31XhbLfjKF01khwzWlvpgBQ5Z8bxW1+TC6nwITlHYFgFY5cPM2BYgf01Cy3f21dc3I/c/S
FbRuiOywcz1LVVizGhVo8zaIPuPAgn7131YQvddEX5OAm+JnPy5LfhY0TFdQ0IbnEWpkBfQM0MA3
OlDezC2j/ElxEFrPiST1z8ApSSHC6ja0lzSw3nnEZviUXNt/tTARMbEJzrJ+3SdTOHNq2ibWRlqa
WYQ7+Ya4W9yPyArpgC3lQCf4JAd8obayxu2P6px952Cafao7XjBAPBw0xSnc1XhrtFbSF3sKPlOl
HIkvM3zONa8O536oDRhdaais4Nq2tAncz39tzl7sXJp9LiL35HiEZSoDWqlY1VI/l/TQ3nDkBn1m
Tl3cRY30GSUKYmjFqRfQsIJkEijk1GGYR2V2E+yS0/VdZ0xbJ2wB8uxgJp+bH5hZnuLOqw0rVrgF
ok7YsmobuBg4F6MCPQ81IEIMxPBpvnx4DfmN9dco12RjUDMQckI6LA6yhh6TVJcs1fSx6mBqLZu6
jnBZGfbiuLSKuTmk70ZATes4bpyEix2QCaVTM3ZTslKuWXzvValt7MVnshEKPSzjN+21k0ZU3EiO
QC9Qk3GLVTmkrOPQ+5yaoE4y+MaUvLxHBVY/Ym5o9da68oEH8vWglIXzX8Oy8ToJC6SjmunJJBjN
ECHyVQmB8n3OieRmp9esrlRiYvGp2TwOqpB4l93r4lSfS/mKJsQCgJL6d8P6I6DJUK6JNnKU8+Kz
tIeL8M7xqhJa7MLqbWbkUHyDssK0r0o3OC/21vHgz21mpzsvOvimv3imand9xGJHpqv7HrW8JgG5
qvB7l+ShX5GJFVNmqFk3nx0C9fKdstrdDdW5v0dyzJ4whCL/ZjWsLlIUTp+OsS3FXgQ8+HG/aG8/
E0SxsI+ED6U47lgO8HeW4nLXx9CtqKrrDxWoK1m+bt+c8AEtzLx5XT0iPXhMg2rMQr5xI9PDBhCc
c0tbZfKOI9DyrJqSInpEMpj1QJMDgfAYafqNPX/w1HLhpCMvww/45lRpGcqbUnEUOy3wVrJJqzKP
rfD6RSL/mxvc7m4ZXFOjPCHZzPjNqsAnND8v3sRrvEw6WzX+Jqg+pbejgv9i6DdemO3ZWhtpTCoW
3ALdrikVfE3LOfyvc0OnSZBrrni3KTUQp5kX4p1GFK0gZC+SBAbAJjuJVdQPORvfGzjaj3mS1LSK
noUZTRAEIeGd/H+Q7J1sOfdugyfbVWvXzO6JXIRlPREQCwospZCoLNgjhLYbryslXMRMvHFjR58C
cVpZABDa5lS2LEpX9qJjhXtjiFSXxtx1QfTdj0U4eh7q+7lXaS/X4fqgYAB6s55RnGO1YtiglSsP
80tX3FBWB4Rai4Pe8Nf+57e8zPhltfKOZD3+Xz11kpM0Um8HMFIDZWLlOzsm4YAH9+uhhwtZ9GLk
LDk0vNzWtwvieIMB+swM/+PNi4MhZNPuBX+/whKI5Kt2SWllJCV27iqNNYzPVlMyxV5Ao3fFzpL7
FE0/Tbm6DcaCYd5DBir/2jsdZG48qz3YnoGYW2QRniheXAXziBSkfeSnkiGsWfI0fyef5IHHSihC
iyk2GOoBT7Q6dKRRjR3+zTEw4miGmmJ7GJLNH1Fl+SohvhzMbpI6ylYCnGRPT6Pzs2Zw7Wag7lnn
e1D2I0BNxsHfPTFYdlzEwQdOQutP36QM3JZJrf2bKkMyHaKrFbKSh22lyVkn8pvUCcokjapkUmMH
z1BRhy3t7SSJucj9P6lIkyuryTG3KJY1Ifn8/n5DDYDu/HmmZqVuD9zHziUo2AAawl2qadhP28pn
qdI1pqMp2osRSrEB6YdpBPnroPkK5vG8TPi0dbF8/GGhVg9F1UvPfB+xh3F5odb4Jrma3zSyiLP8
GWOpymsImQIQhzcW8bX978DeXc7Fp1/QqSkvyuZF6whSSOI0OSkFHPrnr3uJsgHmOZPYFMvznOlL
P7cG2FLAEmnH6sgo3g5RmFthQ/Y9/KtmL5G2HiiwjjOkiXGiuYDYkmNBJRXe79aZXpuAvpxlsP2B
gGtddx9PViTlGP/l+jT/owODMqHKk6Piu8QQ+ePJM3wvp/n4Z/fvoCCt+PMiSOn/PNy65Rou0pdl
V6XlHnjRAUhdikGLn2hp6eUdyskCGPv1DPgmKxvYPPdUxgxwp3DMgllvHxaev4nRy7Jq4B01HKFb
yEUH/mw0doZlygJDTRjapZ42NshrFr/BgvDoDCv7ABJ5IWncmDtkmg55zFqXBHD3qqlMqOm605y8
eS9kSB4CRZ1E3WtGGKTt+xO12J/1bAFnDUeVdHvc7wbkwLYl1tu9u001RZuyoWTrS8sJ9PPyIz0a
XhhiRGbYJ8cvPepBOBgxl+K889o772N/H2Orpy8W7e3Hlr5DRcCrFlX7JUfKySjW2vg4c7g8cU1J
cl1WwhDki8Ix882iDAIrg3cPWqLcFnxTx5vPqAx3fTkoskAaFO6jRAz8HgpKNshABY2QAQBAwaNv
X2HAz8cGEUevYfJUgrOxkK4iJh5bqWM/qt6QIRvleJOrf81Ia/FggQ6/QDFLuSsRbqVAO5A6kojq
e7wO3RFABFy2HvTzrzIrQkfXzJPzDXuwL4LXNeDSuy93FjnMffxe5fnWaioDadZGiL68Rwctg23R
dmbTwIRVMex/djBWzsnYuIFeHfK3V64deF4cMljiBmY6gltx/P4O3bSeYpIpX1KTNm9kv0pnlQoV
rHBWyVPmwV0kBWWPCle3Vzoo/vtILdHqTQVstFtcnG9Rh/H6KfeI6MmS6SMillh2Y3uhWOzDdyNR
ucwqph0L47CbS3yaYkKohKwRK2VW38x+w4bzsJD3UaFCxrt+3Wkx/eiZZmEtT6JBx07UWXm3kwbx
ZXdBV8xj9n5EDlslBf8vgqBhaoBiXZdmITNjlLAb1+pZALrJ0wZqD3qvBxF+pPk+Ec83amCObbVp
5VAoPXiAT2GU0/5ledttC4jA5fUR1IQjKyZuMOCPBZsao4Rx4HVVvxOxhavmOv5TsFyvz4LHu2D5
fWWJX97tEtn8To3axODzO+0rYoqABEyNvuXGKWcML4k11Cuz1phTCLaFTYII+NZBz1u/VjLja0qz
zTwb9qWNlqwzBaKwRKk4vwCxzpA7mzWijvkCKC1vv48BvY9qt0V0jcALPwCpFvPst9qtdWKSzNd8
LxbqUuJv6dmzGqaB2lx8tFvuJXPKP0DCgcywqI/PsJbfn6c7yPmyZHAkj+q3ILY9AAYp5GTJIECn
3P6wwRmP8kHqpSUQDaqpa5BgtUCPyL4pHHL/sDoRfFQnih4ikmN3s9rNsSikicstrS0BGdReCc60
C1XFxN6yKXdZf2LZ8i6v7H3bFwVM1vNCJKFj+H/L/EjGuv9YLD6TGzRmQKtSuC1nMS4AVEHmi6+g
j5VBrJL6Tn0nE9DJaUVvqg9GiVAANl5RxCEP5A46xuZM7X3iYs2WCYgvXbr2kg9sM2iwy1Qq9Rgj
imIcQ21VZUqNQNCnHLSxuoZE0rdyCZBngYS2TNrA/38ctp5vCZFo/NI+gaMPtfbjJaqH1Jz8jIGI
Q2Mcg67hIdZNKTbI+SMA0uZ6ShbDojXLYAG9tbDllkBI7P2H7v/0ga03R/Bv0xzKuTNbGfkCXu8U
mVc2S+rDIrRpmKDIfztwtOEqzT8Xr+A4x09GvlqwfGvcs+BQZ8TtohS7R9Vyoor3gkXoSf5wZM/G
fb5GuRwN/xxmZFJmvBZvqr3qJ27dR2MdIDiJv0NTSq36ODn7iEl3URH8k5QjqPTInctE6y5t0Db7
tKyPcZvnpKGchV1MPVGB4/qsD1+ctcEDpBaUnj7ot3smDn1SAHALufo1jdzJxyyVFH4buwtHEsKD
AeoqwEkVlwh6fEaNYPaF6Bpz3WDHmp6bdmxEIPAw+iqNHoiNJz6Of3GEytWhIFcLWyaBYXWYzBqY
kqUSdINEPCV05ZPXjDoLEwMmWlUk94Y/I5pwIBrL3Pv0IKMA9UW2Il/6D8NY7AE1R6tqhnFr7sWo
BYWnefnBZObCDf5L41qSNsPduJKoe9j9EeJ3KfSoQ+Jn4Vhk+QBNzG5UYPFmH4aj0DR5EYVddzre
8G2lqVOEnCr/rXRGON1YjPztFjQPbt+bHq8p8wATh2o5kaTLPhPdZDRyHLNQgtr4fQOOrGxtRszi
paETKbndiLwYepGM7xkw7KfsgVd7Ma92pdsiM1JMP1VEaHbgbHCH60Nj6CGliaIbe0MdWM32SKuW
RCmnavhM7+rQhUkImGaRBYv31wKnWbmOjDU2jl4vOWHnNT7daCu14FS2iSvQLL81odEvZDdoUxwD
bocKvDIOvtXfqPHsfSFhqhlpjjjdByH941eFWzmvErvQZJl/Ljj/1oEcoEGEuLAeZ4jOZwentq6N
zfcZO1CME3of+j/Ywqpz+uiVT/a5ujnHFAKbdaGfMJYuYDV3bCs+p+JnM0YidsDpE8X9rMY/GQhy
i7byKZfoCkRlKS+CzWKTE8V3Zc/wgPYVoJb8IwtUzzrZiPWizG36TTPURceukRaaE2m6h+Q3gqf8
SU6HwOaltKpcWMqwDQ+ZRTHZOfWTR5mq0Me8l0ksyTWW/Hmkiqjpiu7hQGsY9VNVaQgDbNcrhKNa
PDwyL+Za+8/Veo3WwLdZDbvjU0RN5bg6YaYU/Bdok4bq0PhAiyQa2DPGBm5SoIbAYXnZdn2ZqNgZ
SgupNhRJ+7bks0OiFhBRozKXqN4W0ch5cvjpynbDcl+MqwWPlIryoho8vz/AxMd+6FJu90eOSbar
3/lacQZSQKz50Oak+DRGC19R0EkSVCtXs7oPkW9hUyY4oeTCq8InRx57rhyo1k13zVJRIi+FrJc1
3cH2Kw6g8O0VNYq7lxOG1NKh2QRxiktTn/c5Oh8EV3pWcCs9nB94vLR8mMKELO/UQDHd8+z/CVNt
ZG3Wpe1F7WDDUHgQK9IaeQBi4yZUfD3FMosMkesKH/W5GpBUoalR3Z0CzzmUFwANZyqtwDbPD6Ku
+02phwktBkNVy2aNWaNEmymp+G4RjH+WxTMM9iDZN5gI4ZXadnl3ITk3tqd3Ih7WInOYT6mD1PtO
Bd82D/y+e8zOxSuigQ/vx8+ttqIqpovv9JzB2Sh+4Rjk8RmGRz91fVNAEmOisxDsANrOwFtti81w
sAA8sFiho1vFSAufnCXJM+9XTx7vEUfphi44BYB6k+9zm0M8Rck8osejImnkXRV/vj4Ma5/SIwPG
oqsPglHMzgCLbU+Geml9a4lFIJAEXElSkN6hdQf1Vv3dMdTmfk2a5P7D0aN+1IVXHoZSZt3ydMYR
qvtZ2/KwEoPyf/o7Te8gYlZ+NXdozBmeJpMmfHD4gg8c8CHBkTEF99+Z2itBtRhS5ySWP1lwc5y/
sbQ3cqnUx1dk64Lhz5OPsg69yrPj2bUHZHf7qghsmYCQ3MoMhgPo/dABziP6hZkpTjDk3N10kkmj
Km0oPnV/ZS4ag1Oyn7jMAsd99waBG6KIwZJOQNoCRNKFR+ogHh4l0WS74YlGOg5bQCScUkIridlN
D0tEyGYS/R+qJq548S4I7/B8Tblkw+VtRyE0KGfXPXSHN3H/EMN24DIU1OQmOtDyoOHf8e4Q2Q0m
fQTXh/HWLHn1JRS8jqWt0CcqjDuBo51iY/I9/b5T5YRVRoXsYZckGWYEZGf61gm6vfDyDVsw80gf
H1vA0ppAuDH5kkV4No+KuRvVkl1zsim8m6fF5gyp+TdOFQqdR9YiMCbeZv7kJYQ9GG9vXhNSxbfh
ZRXwLBn3pEt2wwzbjZumtrVNP3o9J+z5fUconzBNbySdkSA9G26OqVaBkJiRZLScCJb7tfVGWwro
WOEy2wB7fG/QMfXk4zkxgsDSSUO/WbQ99jj1mCqkPm7kMvEeEHq1hgk28QSow0loRrwUUgb9g+RH
UGot99yofjvO7DAEjYLmUAkr3D/4VxmDMHMDwEkec6i0aJL8CKNclbb3Zf3CEishQ1IJLg2Y07WY
YySvv7b/bKyZ3tY8PeAiu+/BlCCLTElVK5xoALcL0T/6/mYV2dDmuGABexIx8NqUXzmjXY555zQt
x6QKop62/WHiG5cg5leUmMJxTlU50LUQk3VEfxHYqt2hAPB03wnPopLOaKRlz0oa5Xdc1hZB4EoK
u3c6YOZHotLzAvaR+xMDrBbifyRNe3BQV4SHjz5e6SBMveQoh8T//bEcyxEn+sC71e2LhUvjHQwF
nH0t71qT4NxwjNNWZhb1XygN+UG1PKxZ0kLM9gboj4wu7t6HMxBR7NzNlqgQT253XX0yIRgwzJPz
Po5xYkVTTsZffFaRzvhP6zAUQ3iNPj3K2u4ealwhuWSElqHym8iWEzT58KVM0sxgi5V7aneMIo09
sRrDvc/QhpfPAQqShGTcevSjbzTOap6gg3yHJgJYJkBC4F145pmdE7o96CQU3H1Cb5GZkhPd5ZN9
1aQ3Alhgo7yl/zOUsvPZlGNhF6NDIzo+sBtNi9f+ZdBF0sWGTwWIC3vABmbNabCaQIxZNeHpgdyo
2xv8P2nPpPDFTIK0V9MVk4Sz8fTFd9sKdRkrdkV2aPXYDzJwch+yrxq9Dr3OvxxWVK1WA8bJcMaf
1TjuUHaYetxG0Df25/nyNAWDkU9/WfovkeloxSAQVU3vE+6D0fSmdG5gnm6mpf1iV260I73DlvXW
bBluQg0lgJVt6vFTF7RIMdpzmj7HE1xZ/+R6pCQpgSPiHsJNxWmeBr19urwwipU0BmcE0R8JE0wE
RlYH1LePnako1Qb7QDywGTy5xW0jw0kcGD30mVndgVnHR4qhBDUxiN9OIccQCg1jsMXPINIBD+U/
SoZFwe6LIY+BqcwSxCV1x9wAYJvhAr3MyMbe73IyNc5djjXxpFSZe0SPuptV6vOJQjS9xjH/ZW8m
8nu8ZTCDDHuWyoTzKguRidVUnYaOQi7D63Hjzs/KouCwm5hNv1CfugHRIfvb1FU78TzM20wWctjp
sw6Cpup8MXkCxEEJuExcjAc/KVQa+5IcySw5PfgiCyv89I/pcig3XIWT5DUERYzaLOpfwiDygpyo
/y9Rymbf00NoQDe9UuEYEbV14MwOqjfrr+Sr+JBttwzd6AY/VJF0JdtEwV6ET3VeZM6rscMXUp0f
33xArdZnYfzbe5ak182f8tYmV+Ih2tfPvX3Ytfwh4HtuFTgKIXHLGM9V2G7MlbB/8owlK/anWvTr
3rm688vdeCe/YsXXfW+EYkQ0LpSotDvBpszzPtS1UD4RbyPBPn7Gc1noSPpGAkN/2hPy0ZG7yyRS
giJbXw5XB1CEsTKLrAWBk4OK38ktCw/CUWNpWy0bUI2SIW5NoJZBaXiOw8tdV5M1RN+qCOWDm6RC
XGZ2aUc1T6y6NNo/Vd9OFPrY1kBzzbSYJExXKsQ5b/PvuTCh6em1qgxTfy3C49e7TP30/+rVudOo
u0dIIDJNNi8a1lgfpMvrS4MJbk9aUxW1syqZRLXyYpFJSpern+M04kbaY1vBlEusXi5v9bJQDKXf
6Re4zjABlGOr6wKkHQBOPwHqDqmU11E+GqPVqzLvBU4vuUwkup5GyME+p5NVqnYtchFZ5HL1Rc3z
axDQqI3JonM5mEAvXU8/XFlJUNAjMEkVZEaH/+0a+HQkFRNgQan5gMHdP4SBnGCQczZ6yCdUDt0j
UP82SNh9R5PkxNkz+6T1Udr7WMsh+j09k1iN85bKBhw+eLjN+Dv1wdehcqWWEPU4vhtTtvLNq0S0
lgTw0DfkXXg6Ls2LnV8d9O8J+dBogzItNx8N1ABPRLtmntAqKDLiYw86M7ZoJJZoprR7vX2+KLIT
rKSd6mBSXLYLabitjE7oTNVRmeFN9A/50WUFkUGdOeHKPrTUJwNJhl5YnXmF8bY/manilr3+/KTI
pwvsOTb77GTCnOcdq0mh+Wg98T9OGlnlYldJd4mamAM3J7DDm5WaCtlV4WIDZj6uNvQ27F8EIZ2V
a16XVPY9YrgTEvzqEJMLIg9VBDLy7q6CKvqezYT/4h2mcUgSVhA0GzXt2vaCQiBomuMLGtKdS2sc
ot9zvDvVB7sAYXFVALPq2j8X+FLjHNjL5VmdUAcoICW38kruCooePcfrRQ6pldp/FdG7M4pzhdFX
SHgV5NuJLTfY1xDcrsdIs3QOV0n9kM/yA6TICaa6GZWB5+5MGR8l9pmbx19ijW3GLDbxakZ42WzM
glxlMcryVvuVevPN/0XaE8BLBtyu2psxYOfzNFryxV5ytd9IfE3dtq8t2kR8pU1b1VmBkrcyf/nr
4HFg2tl+hAK/cDXmUYKzHTRz7q3nmexoPR1p8JKHjxdZlfE+yPWPFpB3qstcXs6SrFS3gkRW6kKt
Z3dqnz0rXUFDIVMnDeADZlrHgoHYGjieM4Ah33h5b4nabP6kLuCxuxVzSPVa6aaWdR4Tx12FzB1j
Y16xgopvHF3/hMS7QiP0BMEsZOYG8gHNngMXWQeptJXdYWMR0VCb92A5kNB65gF+fKnlijRnSka4
3Bld+IUBniwMWdaMf3NnKtFlhjYejdGdfk17Awzl8ZMBe50bw/Bl0hNDHlcHzSdT3fnKQVY6aCMR
SdfK3oo+s1AGc6iy4J9OlkpLPiqSARcHntO0Sac1VYynpJp661vyzn6NP1s2yI38VAyPVTSoy2ZT
Iw874wcBCiCbrqko49J3j+iInki2KJ4cEYF368FDiNC9zUbjrezULP5zSJYa9TFSlzMTdtaWBA0f
mU2XETr6l7OO6Qg+u+CwfkJ0uZiJiHfqeQ4D/U3xKGOurs409BTkDhG1byqb2tKErQjOl67cHmFN
NdW2TZUgFG77YR1Tt30X5JIgDO1Gfs6SQn5bwxx9JJc3+0aZLD4dVuigDBBT7MKjHL+OFKpE0Sk+
qLOvt9ELLqTOKObS2az10eUQz1FbLaIiAjAH7MMJDk3VjCwRe5zSZ7NlJ02rnWHFgpRJfGm9StTd
g9399yRGK8SmC/W9HW4a0TbxpsE7jEqX+TV0QQwkdaNMJ+pq2SmAyqb1mNZnbc1R1HDdl4mhJLap
7QIybj7BcBR5mjYdEK1rwXeC+CndNDtdfQSftYVgyc5dfMBtlA1axmyV52OEt98/RtV+KPGCCXDP
J5ts94R7K8RSPZPYCD39Wjk9uPjxiR4hu8IFgeLAyftDga8Wf5JA5P3dgTT7Ml1pUG/um3e6dDaB
TSG2ixWND4mIKXhhgA+cATS/mfJ+uQGw47XFFJtYdc5oigkb+lfSmEkCbiVAx0OPoy9CR53Ec79D
UHqI/n37TQulYxzN8C26NNKmQZEdkB0iN8lstpkzwX/aHAWGpiiViPskVZDnkSM6b8LpeXWgw5Ot
Tv1OBLBO2AwkD+hWJbc16BplCTa+F9HB42S3194lhSaM0zO/XrdF5EmlK5OCBgzKI1z/x1Tf5O36
nEsSKKjD1b9UWk1a0l98eOFvbwJpT+UwBRuz4wngt1xQg/Zruk4pbKoHLJGzq+eNYQG/YexYMMtn
3h4Id3BpkXJh/IqWpO4UbqJXawxL/h1TH09ZtQki8ImljfbkPI8hWka+yGLY+JtfK/EhpP8MJoGa
3hOmlxdMsyC0Vq0wamNP4pAd4t3R5HNOnteLfEo6vO1JPh6kYjyXEicOIYUqKvk54kZr2GYUjDqr
Lm2bx0Ob2nKkLWxFMoyoM/vwlYvuQv+uLmlA6r29iMHiwyWU3mDkZwEuSjw3++TqpWDdvYpnWnV9
ptYbPc7EUQKBHP56aWMuTH8TAJ/aq+yCE9LQZcosoTcEkP07XApN2VeChnVSMo7i8QWF1lPkqY3O
5v5voQjeExfRSPNjORpkzz50ZXmvKjyntn3uHR3PLnqtRCvXSDYQMOtQQNUn5phk4KIOeS5xv9D/
F4R9Ah4mrv4Q7NZ2k1+i/PQflW84j/3ZpI/nCLiySjzvsWs8OqIewVbXiQvV4MsQmzlGKZ0NSZD6
9WS9OPDckrWBP2bhD+VdHq7kXnD4bcM7Chr4tpJfFdMIxijIyJrW6YRrNiSCP1P/507IukZIty/S
tTeI1mQKWXUFHpJlnPxM9BhPFR5b6C6C5h98Qi9DUh8iIbbgFLWWjjyh0BA7EcMfpoSXa3/zjZHF
qyQtWb1QMuAsK7oCEQCpBl9gzdTYd6Mzrd690Zga+z1sO4aanw8/S4RisZq12NMJz1CA//BvFyK2
4AbNIWsNxIG95qKI+xmfD1UWFfS8p3zyiTym2bdMI5GRPux1H0qZWn3bBZlJ5p6uS4NaMRIcDe/r
5FfylHm+mRbpd3gPGTFzUfFuOkkgMvd0TwFYThEvv/rrFLUCYp1YiAJtjzG4QZRzDncenUu7B9V9
hJ0osdEcrxmE9NjQNrNzIk9MrWiMRCM8oIRRR5wv4Ddu3ImEqfBM4N+Wi9H58QP2LkQ8Pfm7JI4V
tQyIJYZhrDJh56Lmx01ZeJRja3nY1IsNWgOaktM/b16UJQhCnG6sSZqaAhGfHVNqKeU0hIF9D4qQ
LcChr7KOOFkZmuqT608gwj9N0ZQ1A/lUe40MPn+8aNBCnVJsBE3q2Su0pony7cT6pWjsUYYSViz7
rNp589g4HOvT35jh6+b7qYve+/IuVzIJP7ss6ZeF7gMnf0kA80b0yXNE4FMwkAUGEThk4MDOLjfi
0wpvSk45HLKYoVhWgZXlrTzGTiaYupI05rNq7R79kvW3r954pZGqPHUWNOQySnHx3FJaRVYaFNNN
uMPTFJYj3485343U8dyJjTSnrXAv80Zxo6FhgkdO7xeAWBvo8nQWvUAbTt1W6bawhx0wGpbOR7r3
xIT7EYqu9QmvCAGO32jYqiHwZq9xsqfXnnDjpDrpAeu8XOTP9iotUlFKRL80QD0eN5wbmBXoVE08
hHFLJ1vJz4KkeFC59Hu+GuA8PRkgbkHfavaw7LamWy6ZFQkkgZ9uyRFVI0SvJRipANlcmKJRwRCY
9XFyh/3neLO2Rc/kGWHKrabytHbMCSpt5CUsjzZ/ph6AwiqKZbvjVNMbyTaqCPoNfosrPqGCaXIe
U+gYwckcOYO6bTE+Fd3nF0D+vwJ4uLvXG11nA7/GStwZ0+g1BNsCrfjih9tdKRKJBcfOCuoxxVaj
9CYCsSVEqTyWheo8UoF81Gwe5dPy8ANjRwprUF4scpETf5jO6Lhorsrd16+9JV/H/0TMnQzSRA79
xu2FvfbVTa/a0lZK/YyDnA+bEOUJl/SgXVugATiLkffrr+WRlQop+nFyBvYcecn/0+YeaQIlk6me
+1Xita4nBLG8c/nfXxI1PeFkvWeOAJMDDr3IdNhwtjHzE+R8hCAF4zlV0LI8vJ5K2gxtSyoFG4op
OKAU2WVNj3T/NegbPR6P/j9rZ53qFEKg9XmSU1kZZAT4DwwL5h8srCpEPpVb2TZnxLZY9dkZBegK
A/iaNU2kzsLlpLsuqcVAOygmfp1wpP6g3xRNFMwObpVc7jcprhlXBTNDPo+A6EZTQvcOZr/TPeVy
d759SN9nBZGVaS7WUvBi/bg0QW9YTaGI1q7SamumL9vYWYY/+sPHUCeyB5JZyxrvnn0f/RPNmtlE
duLgqXgewM+FCXuQXaL+uvfn+tcV8cQs7DpbEU4K2VZEmUfz8CZsit8xv10M1ioM2uKmM0kwOMyd
/EcUAuLBu8b7iVTqSfEGilGJZ6X8MG8J9ncFsOWoRoKHTbItLnKGTGI9a9h25doUfvUg+QMbe2LA
BD4U5OFtYpQlGrE9MLVA5xrlPNqS0pPqBDB9O3nnSQXDIDrXDedJ9vXVT7F4I3AtZQLv8LzWxNyN
9UDPfEKPkF/3IbWW+4SBRP33XTegb11UeOtUCqsAyCohHSxCyM2qNht77Wl1qiQDSFx/dwBq94mz
u14isGcwm3LXSlIKIengWyoeFh1mZ9wnloCAIxqPSLbQAllJ7KwBUbJNKzFWTkMYMG1E++P9T/kP
Spo8xGuwCRO5PPndSKd2S1IfaqCtmEh1e9y6tWoPo98a5e++UdFsM+u7/dXXJ7iVpdxXJsSa1Yc3
NtttXpl+dBqIK+WXdEdCwovi0QXmJuBltO3InX2WWOJw7Zw9a4K6J5mQrLMNA6VtwvYrkhbI3WcL
HYdFgYYbSZTqkTgfVBX42iUpv3uWuWH9OVH3I3ipGRYbuyU8eLrm52kqb3zFiMC4JYfFJVsI6Gwe
olPzJiDscOWum+iWKbbt5KJQdFk+yhxiKwgz8145aEWma1JDDBnEZpjn+oaCYBG0tRtedgNquYhX
mKNmgOGNbFzsF71uu3S0OxTmY+981pUpvfyPkasA0RcJPFs07BxrEWA/j6fu+xl6EyJkmVGTdSPj
cmtNz7kYwhD0zIQf9eeP4QPJDvHjVVcsbowpkkqO4+nWUvWaq6ixPYyNcIbQDGgU6tuZ5xBrT/Ry
7C8zoCLs0I0ksr8e82OPV8PKcYtyJia9UDbwbdegBDdan/N5CBFXZjBbR/nbW5WKH2GqM2tEA3w8
kuJ3Ofpp/9QUTYSAdjwMLYPswOMhmUNq8GicTBxqPdpz0O+mveD6yka2U7+EJDEmYS7M6Aezxwje
wiKNqgML4l039Vno0bP+WAxl/Wb1jfuYEBnS4GS+uCTh7nZW3C4AOBJvzlpeEWDAE2tfoE9oKl8X
qVJBqqdIiRG0bK37/1n0OD1hAGWZT7zjN4+VH0v1Qzyi9BSjo5WLw3OudpZkbHr0JkwVR/7iCHgM
m6WVrVQQrMJocR2IUKJdpGlYt8Hy9TMZAkpEl7vmsBD+L9bkyKItD/sfURS9eyKqozi11L6FJEeO
4d7ausUglMkimK+ko//3qKd5uWYz52MkKueCqAip0A19rWrP3gby1TuuDqsNodQxaq+KbnCwvH2k
JgLjI+e9UDSCsL/O3UH9KmBPYTnVewZ8bBIyeFMTnGU7umFCFjBC0V8Lirzx13MqNirQqvmpPwFi
A086sTNN7WLgZ07qASvXZeIjE58vU4ZraivUlbq3wa98IdtrKRpF8Gx7deTp6Soxg9eZTi818nur
DPi53vdkO65V5UKOAIFgAar2cjCdMu7CVvW8XVHyHcO7aIgIP9EMD4EV9T6sfoM1HDVCnOOe2mg+
IECWegJaWyGrROOww3eCgtB3sFHSFcs7NICbs36b933cwmqND8L4czS+Lvev7rGl3OjLuJhoexFl
YEEaQlro78B0E6ySctlEVo1Bp2iU+hbaSPA7byvjZlUXLh7aLnzHvdUOvPugRc3Dv1UJQSuAXT5o
A5OJmxMBcYumE/2gDasV0/gz0M4yeF9Z+We/10BFbsLEyaqwNnL1J0RQUU83K3eT+B6FhT6q/r56
RYGJJiOnFySX7f0/63dxeJEE1+Oxzb5xARgjjDaFSmyRDKjHxTsndcV8bVQ+A16MjHx7BhMhAW3Z
DN/KOkVBhxkaIIK87EnEAL7cqydIOrP9Go3GmyBtjJYxDfzHZoTNVERNdYByLxOaff3aB6U0sW/t
T2OI2T4rWp1adAtxSri0FJAx8X89q9SXeS9h/Dt53X5av9AOmMSoRH+oHu8MYDL7udYSyRZfPoc6
trOmTIw/YMsF22VAWzjOhqvS9TXgRIGuFlq3dS0jRnXtb4dBGhoKyQ7S0YvjwxZVRRztUuWG4V/n
rLB1q/iv184kn2tvgFOrcQBZpKfq2e3tYzzKkjZYsULmzYqIjoNIeeB8RFZ43QSUyg/VmzGJUHaS
Zqp53SzSLsL9AhzvRnRL+15kqPjMdGnJwZTZXSqY2HJc05IsOTXjvOeF/Hbvab1xnZNijHmCnWob
K8GBNhEHnLCmIFnCYFr7HJ6tOIcetW604fcMgH7NQ2fXUL05X/QbDBija9TDsRjo7ga+qXJCByN6
FBj29mVlRKe2/ngYP5VhNfeVxUGx1v/r7muLf6fYUuscEEyO3rH+d/cpeoLLxafl71mkFXk0RbDJ
tq3X6OmLURstFqMGJoFxEM5tHpB68L5HKHEsmPYR54g+KJgpqFqhLnor247Xr6xU8NAkWwFYv6QZ
8rOHJmNmtA+vYQvavf6/tHG5CVdc0YZC55x5gTHu8b3sg5MbCeJZvvf2OaGThPoMz9cLKVr7oOv8
ts0R7FkpUZntwvEmx4jszIvZfQmUH8D1xmwcdAFzNwVmCNw0VMgICV3+99hS52ZkRBMHYgaPF4LB
kQS5kyMGIGh+feVTvO71ob+5gLgxHtC1NIoE8gjzncsc9/JsiZRMWi/BqvLQNZ/jPf4P6nbl3zOu
+zlKVP0w/yio7tE8jnX0MbTrqWuOWNp4WN25jkA/V9k1FKVAkAeiK3XlNimqVL/to5bjRYOJYkiG
/nsRqz59DcehfdnhLCIuZoBzE7MJCKJgaDfdPhv4EXZRxdG7wwETRYdNOUGNFoRl2ILYInzJQRhE
MHAnlBXsPxKbRFJKh1uOPX8rPCPLdhDJ6G0LLAwEZFGASlWv0BfUQAD7nIwpjmvk7E1LtpacDmd5
6UWlOnwZc0gvrJ3WYKz+eFuXQNRZ09fPcvJ3HgR6XrywbjULbfoPegimikZovo6H7BiI58nCYOhZ
71n6ud3lzGpvITejCEvq1s3v0VOTBg6+//4XVB+Eq0jZD/un717YhbwdsPhKoOhwNPTUOb+SPtHc
Wxxzc+l7cVmBwWmeAZPdmSk5QUzJI42KU7pnFBC0Hr3mzJil4WitRvr+npVvKGGPXrdoMGmy72Di
+IuLqi+ZQQIf5H0R6Bq/Ww7m3V8vq++L/lpRpbmCT9pRTltGZz2/B78f0AkHSv1EQYEYnDTX0znH
0XysP3UfR+THhpTZmVJak7IkIGMyBhXd/0xQ94MblZfLDGsjJP9nj9ZeWIsIsjjA77SeKjJAIkqk
QPrBBtgZjOWzCokoLUThdXdjBU1qPOgcH4VksRlzrrf9ARp3zeIjhsi3JhPRunha5CJNwoHupCaq
6WGQtYkHLwMPy0AOjxyY1Pi9aCtveRNcWvnPv7Fj5PYULj3bAhezdiluh8o0Blh8N2IZt+qnpzhp
v+P5TBZ+TxNRmEFg8jdbkdlM8lqDSUhBYq2xhEzFV43CS5+2laTFwzSI4K8bVH+62efYECau/CRv
+bboIhpPYf3GWK0No3lqqrYQt2wmhgANQPMPJxumG7JLHtVP3tIldMbkga9z+W4l0+zc1TBkfN5Y
NFTzp4n1WKkz7QC+goYB91xhsnz44Wog/y3d9XOJXhXJ9mPcmLrVQbSs82VtlnP041oo8YOPgNjy
5Ji1oHWB4e9JlXBQVsIpYShVcQSghIl8/CPMsZbTLTooj4Z/wkVE2xKXqiH6kK1M/AVl5o2moFYp
YeD7Xs6s/BA04ESq+0zXqkHT3xBBRd41FDExKM4tr1Usf3pAx24XO9ejnrN1D34nAiVzuJnpdXgL
Jnr2YoLkhXrJ6EpsO34Zf4NwtYtfLGZ1cTBIEBfspGQCDG/WcfEVpkNZWILJqkFRNRZIIMK7t6z0
HaUrJ8n7iUAahYIOPtt+bMWcc0eFyRoCZpyZz2TQwMaszxMf07mC5N+ul6/sNutiP0JVJiMr2pZM
Ni8aZnFvVvCqC1O1qVueOulFhpxMRa0d2qZGlFEAV1zHOwOmaNcD5Arykq4MCRQyYxylwjimCcDJ
0DoQPcyL+LflxqbZAu+ABP16Whe+rHSMC20zYl1h/r6UdGfVW48vvmroNEp5Djpxfr+L30k0FO7W
sZc3t5n8woRahxGu9deeCnwWuWlbzyKeMp7kqrDxR7Dol9zCcBL/3GdLslIr7jNMtNMQULM7j2J2
36cfT/PWDiJ+07mDjBEA7U6hIc66oTi/B+xEru4NP8UkW7VhqON7gGtiIlVd0hlSuiHPpiqllxUT
rCMu9q7ggTrzMQrFSx7flsTSubzaK83qvFc5iNd8UgNsosXvgrJlkDO1n7xTCzGO666VVAhVuEJL
oj/vcf7a4UV44Tfx3bdVOsrKQkSdGXVZ97cRhQIEQhX3RN6nhir9o4gIqzPItZpbBtjXrfXH5bNL
WvGkSo9/QCXrmCZLcAbb5NdjjxgJNQ5xl1kJ+PXdXYAzHMkCU2ArdmDhTmw4mfNgAkCw6NB3i8x8
FmCXLD1hHjd12wfi1rz5DzM3yI4WURccEg6tpmROcLQhIEDlhvZqW1BmiOQALOMcWZbqGZun23KL
z/8dUMt+mcLLzXJHOMRNgAZNtzXK6SoOMznw8992246KRWN9NGto9sYXP9gT0PyM1w5YpmHVe75L
IiaOHw7jS9giVLz8tUdo8OdZ6VG/wnPiRA1Xq0avl1BJZ3FYRgkBNVPPxLInDXAYPJIGzUz0xN86
CjUERbI6v6/a4qNXNhdOPSDBkjrgm51S02xeNM3Q94CxTGnuNxYqYb8T0iMbhvk9T7qoEQi676qr
mSzQGDRb34kfbl+H1y380nPs2gu2koG07pqrA1y4X7CKEm4RtghLcUKDFYHaYslnnOfNKgvXbNV4
Fe20jjYu5LfPb7U+0iZZpvXnfApAk8UuBTswwcGS2QNo3Wh3FaYYNPEFyitOTmO0YG7mXSVqpHu3
0OyCpwK5PIzNYKwe6b46pvm0gc/qMp6BkQ4ggaQ6IVUlFX5FpFYnaS/PXmGTxRfDu/KxKquSKcwl
ylF99ZAhSRaIJXZK5HRUMUUea9JyJIBnKC59SIRh3/L4gLHlWKqFvhnFyFnTnSx4oJ1TjS/fOQYy
J5G0BQT0VT31t/QqrnwGD/najXjOIq3XTrwmIp7FiMIrd3F+KppNh1cvS1koFvav/ZEtSRq/A/DN
RnuI8xmmRBK4JtpkJgKAE+xhJRzx8NTZeXlb4Tmv5VcGKxos8rlmlFgRogtuCDlZw38+zATnkkQJ
1UTOkOcE1dXjMOdVdFkk5x0QH6u3Sy1SV/KF+amkZJfGbYWFqlkVVEFRySD/lLl245fXS/0A73so
+JOc37p2UkHlNwR7K8Yd9l3wh2xzoa6JZuS6uXybRwgenU9Tfo9PDAYisV7ScuiRcthD4r7miUwY
PEpmEQLNUM9BWMcnWlobQKFMKXBnFAUX+PgBpZn4lCYjTev5MnH+4olpvpC6KM2P0aaWSJTypN+z
5ua327H3BHcxVwAEFL3S0Df3kPCKwBJZJYZ57Ha8c748BUgC3n7U2mkLtAUzL3MnAfvedOoAxc2T
78hJzIXperGEbKgu5O2CWObW6V0pUKjRZytN7QDYcei+A2vGUW58Lk0q8NLOsDCWW6Zlp/OetNq2
vS/ywtLwMN/iV3xvXq53gRS63oyQsFKKzUx9rWtocqz68BD4U5mXnqx4FhFDC8Sl8detrrXrhuh9
oAqnuimQkIa17E4097fajUP1/8YbWyctHsRYZq78VBQgpokGVxZU1gxFelRURV18sAb/mkkxhXVU
sEiUtGxqIK8zMxzxbifWKWwWW4yn+gXsZMOdH3kzlBstPsy411rKH6rsOWLmPTB/SHh1COwv7LfY
X4ptANd6PKHufBElWR/VfSZVnsCFQednbxM35CubpK0x13z7CYtg7FqIojOlD8hPtOnfpAMgIyR2
LhGDc//EvA5X8cZyonhENVMCyjsmLlZRETpKzhWNn88n9kML+xQjwZ7/c7qb2d+eWPgiaP0q3Ku8
rEuOpM07lQsfPsb07spzXnNB9ipjDo2GpgaIxzZlWcvVtSiFkQ6zG94x51e42jGTfMc6odwhFF3B
tvFMlDalaYFTI3xber/07V+jEnbxS4Kp4Eww+X3dbMlle/eh27suI8eE8SdVorjt+akeEu6WpYTa
Q817zpQIERTQo14S3vp2ehNMkcMRuM+PRwlzZ8cq6lGsACcpUuUekp+qMNxamFjxuXz9ybpiTMn7
vqtRPB3FnQL79TltuvLDrWuaa3AbgE4cfBp9WnsLsRYqaho7EGyBo48SENA8A5tVa5BDJXcdzr99
+LsZxYGJBfXsVqQOWdTwFybVrr5+ZfE7P53wBAyRbp+4ueQ5g+idWesguQy3+dvrPBsiRkpH0Dh8
VoNb/2X/5BPVB2ALvinxOsPvceF79khNqXFmeYh+skhT6Ohm2uwrmmFXxd9/fZraDrOly8Gd2LDq
Wd6U1ML6Q4Sv505Jdc4tALPRaU9wUAxFxj5Wo5VOfOT2g1XOGJw47cx0r1dJ6KB4/NfDjDaMYZ4l
VFjSwylQiTiYGKeU6SRqPdweQbDyN8ql9pgYilUo5VDtqHcEfusD7BJPQA3Oi4qOGqrLQ3AG8GS0
SKxA2s4Z1wNvVa9hfrDy8c8vHo/L27T3Uk7Sl3RF/wDfX8B/8WeOqjF9sspRCOZwOQoE9kVmWVIy
lk+vsflnlx8E9CH9XKtStRiwYMqfq5Ip2c0P/tmDjz2hir08GlgM4GZH05F6D21Q6LfO2cpttGzh
wuCdOOp/V7LRrfx/m8tJJLpC19znUPj6vt2jNA+kXfGU+TxVQA3mh4brrmI6XItiwv0qUxdX0twj
/iti5Bc/KeJG00l5JvU6gsOumtVGWNZ1hksnW4IoP6CKFaB/xHd7pD/kutl7C5fmAvGdmIgvKZw0
AGbfQ06pYaH2sRA0XbT7+vpAZ++6dExn+Iz/SZ0i3wAjJmbLpVvzUNFEC6Yukgj2KF4ZfwIUwvXf
QBIXrj5tjQWXNAZZUnapQuhz1y6icPcsH34AKpZ8IFskKRULLZDTMc9574Eom1jiAjB5TsNqlOyl
vnIHgWtXpJtN08jpq2lNUjo/SQk644spiDRkWF12BZPS7iZqvsxgZYwLC9a3JAsH+FjNEXH53fHK
KhrTmE6BcMFGOu3bmefxoChXBqSIJKSx0d/lhJ7Mf5a8Et0AeKkdfUwN5/cWVevQtTotP3hVP+7R
aSo1bIgSPYE2dXKhN/kdLxTYerc4sObaK53WuX5+J6PkyuKYzQ4EP5GSD2p2m+nPSW0rRtHQxsdd
zp2/ig6PCBZDVQMXuth4j2Hij3voqH8VGMQSXImun38DjBXRyn0hhblNgKswQc7s8bslpW+0pnVT
VYeqkz5C+j0rYsH5BXKcMSctjpUdElBOztokb/m94gYt3BhR41bCju7G8ToUgHLprXeZIWb1niWl
SYZkVHVLngiwCCxFswy2fyEwGF2rmVtK8CGVv1+Kh9hPNiAXS7Skz3MBm4sfys37linWSg/DO4+I
MxuuS4EsP7uMrmbkXcgVLhlmCp38zgptPIUpmh4eOiHw7OyLRe0ygGorFrCWtiaQEKMKPdPRCjyY
nk46ejgUGahLL09kkjjpDlFytdxaYfsCRgwmMVbGhqU9eW1L4MQjSzQZTiamvAtqtoU0K4GuHU8H
Ae//Rdxh1QtiMoFCmosDUmu2BW6NaH5v6D3ybzSNocsN5HITREuT5fSbDhUxfuLgaiZyh2FcXahg
Z/sbskctJ7qso3RtQgjOSCeROn+LuZyH352sw7N7oTmvK58BrDMP8cHA/IK8QajzQJjgXCk6j+Ww
Y798L8Di6m+VQ60kZwoM37u7tT2lr8dwR2uqggp/yqi6Jw/b++bKFJha40mmTFAhc2iAlLXETOrD
IPm65B4kXJbEJRLgfu5yz20ysJL0j/MfXNiXoWK9OtCjzFAnaOsSvFXgZAfERlXbDwTkPI2JhAd+
qei3PYbWd6Ts6yW6AJ5gmdDEHoO07RDfIBy/xL+JM4itsJ9ic8XS1rJH/fEbwpMvovW7bW6dBD6D
sHncFT/z1FHQWjwAtaCeDfY+VvTp5GEX/QSck1GGiL1kFkmedk8p5Ju1/GZafllTOwf+WXG/rNyp
DdzwR4vD5i4g9t9K8igaG67TkZ8iQNcFP9aJg4GygB+L7KWXxNXmr2lhmatS9GFcRTCw2OEj21vJ
vgq05IN0EWDiQaN4/+L8qO+s+Bi3be+WY3wSJmRV570QsL0DUpi+gvrM+El4COBTP2wfnJSgwIxK
D6Gm+9ErZlLjQewehYkNIjW28Wg6sUsCozyclvOOGq0HQLPc5AVkWS5KjMBLZGbW6ZPf7LDbezmu
wSU6wrLia9fqMw996vKW5iD97VOt4D9lGfyd05mc1ennINUGitva82FqNhfWJnTfxDjQMeYUzL4k
hfWE2E+u8aWlAqG4Rk02Y6bTTzLY1VlbV3kqWZtQsvXuPHiTPZdcubgC8sKXaHbhfboQgBamU3B4
8++DaxLPKFXSMTzTWjxbx/jiltGDDcsYTTs4SlFqwyVtK/aNVJ97HIePRFxHckeQoF9ZCIbBOJPA
L9w8QS3uhsfUP2LsdEs6fRXYhpsmu4qrcXtuNIFdV2y9wH9CnR0EneEH5w0Bvp7diTEUTqBlzrwN
8FELpOE2rcgy/4XGuPtiO4NAnPxUgxEdFRh1rgfnCRCYEqpwLpvAzIbtAK94epAykBOxXE2HkXtR
eKu0FJYXO4t28Ra7G4pUgmtjNGC9R1IQPSHKs6eLHTvsACKzxW9snRarefcVf9W2u87wR2NSfBle
MKE3LZJBw1qcJYMvh7OR2B5IVLR32dlQW25hJad/mAzJznE9Zwu27kNqzVFndYkSROoLQJ7vDJPT
SJr2V3FhbuERnZgtidIcNrFZIQHwS7Gk5KxkWI1ZgpL33BYH0KQ5/CYBmRvE5eIHSyKmqL5DFDIE
Xrrs9W4Pnwn89v4B+vXd8QGEfK44zonaj1KHFeZi5xJPyp7Xt6p4EooLnnuDENGqWsHKiEUm6yk5
TpWpEIRdkI0HCxdSEqzWGnnonxA1OkCHHFawOq87F34YBwwZ1xBQ/LswZP2fc5xLy+dS1e+rAGi/
te1yB5u7SZPic2U1APCpHiKEwjeRjmRb5wio3KqNaVvAtUpyYoS9lbc+pv0NHnBdptXFlnWO3zbR
NZUdpuhELVsDmJ/xXKQOilCMB5xrrnR3eW35AuQafU0qfeQkrvKzIXAO7unQzL3sWa8NKFM8UCiA
2cK/fl/L4mTvSwvI+CeMF1WfxdFQAuBaAwjOE9O53MjBxac5rpiT1kD1jKCZlLflQYbn2EoDCb30
nyN1CtFWUWTGAmyhpE4CpY+FHTNaHFoNd+5ob/ITzgIc01IoMu9w1Jwbp3Qx7VCZx0HtWMGRp/b3
xpScaERxRBxZIEsT1VVQHckQGROQs39CiG7uRu6f/Ld6cMKDpvzcBxaLPqq2MoSqhPSkovQDrS6W
zaYKb3XZ39RZUimbzbOiSuEtcoCyu+OQEnil4LHeXCh7goWndsHxwobVzKd/+d7RGB+0vcw+Q6fU
DkbufFCsQJilHcXHIpugYszH0M6pIzA9lBcbs/OUzYAkXAE3jeIGSHUT2z8s95UpztxC1pZlUK1S
tg1cj6EkFbBaTAC+PRcTytZnXvtuxbTUTH3Fk9PThY7uCYQdEzBeSj6wRWyAoDHZNFXoivTAspIn
zFw0x20T8YQSUgQSDGXlE6u6w4EfEFhQ81QIOdPFCVTtEG6ZgSa7tEzr1mau6insTB7j7IbtVxGJ
iSy6x+HVTXVexoq6lSy5EjcTypjlDdYepTDfA/HuSOQ0FGoxPiNVa8bwSlAcuOz7YUddO/SslnoK
Dbq0ctdnCu9YRm7CSLsqxMrdmOD9l2v2D5vrLXSGTTbuJZPKArmbXzxHMGZoespXieIYFpQNRujO
HsAtWvLW7ae8dum0K6rSc4QHU5ftGmIZZXzd6LxbjKXnN4/LqzXH8c0sazvIPhdywYZe2hOqQAlI
yP9ho7KzY25wXnn+N2LYfB15ATF8+ULVgoxStGyr7gxfByi4HCJutwU76iWzB3rRG0IchmiL9O4n
T+1NVa+/tXg7weTFBXZgHzzTILTq+R3s8ip7TTFN+YoHrG8HKL0uycXJ+wcCDj6kFjUWHpnm8LTp
aYcbpHOWtg5axFPqMBewtI53jxuXcfEDGkhA4I6+42/X5336pCou6M2kmSSHbSGccuk40qVKzF5I
6DypuBHwLCUUxIUiZBB+aymDRpUyu5BOMjLgitcUdBWgqlStBzrfaMMTMrqsJ0WrwAigLpl6nrvm
Bm6X79hB91qbq6cd/SwLjaF+LRGdwFvb13xYEKmCjvVsTHiEtchXv0dDHhn4OGiaVUci/PGJSidI
cXBFoh5stsTa3iEXxFkjigtN6U6kvjjAoeH7Yuf1pLSvFtSTuEIdmt166zUa9mCkZOikIovKm2um
sR6KKMPIVwazPppUadkjPjIMTMxEWNIjQDyZvKRF2gaKgRnHsCkhQGN6eK6fBo4I9gsTrUrHFPcz
TSH2ARDxJNkq0FYx1dJiqp4mnkWLBHrk50GN+TMe5iQdnxVF9aP3kGVfXJbycP8nFOjTqonLR6u7
khMXVzG7W8Z3YD//rwFyN1NgFdeMqjqINsF2CC7+mN50QcZxTC+PbJo0XTfkCUyiKWEXagqwfiwo
Qqp+2tOTW1f+UTqx7nbJfBT+fzHm4BHgAA55s4IjF5Jte2bYR6EnqnhQFD6lkkAcpjl44mX6mBT8
uJ4clGuKVPyCpL8draJkmYCxYhQWvpKzB6sL0bFnaqMXKVDVv4nBsBHJvcqrBmkMwXPT54cVdRYw
yzsOOfeArBFInmOIYFSyvFVH/bPqlbLoN3y0KI39UfDyJjpBv2jwaBNGbB63telPANipKCvdnD/D
UmIOs7Qg/AMbzbLx4l77qBFz86T38W0stLb0aUhFb3yNiyfb4vkNgLTWmqGVXZ1PtReT0LWnADLA
ifhou16Qj6Ftq4K0ZmP5Jpr5sbHG2+y2DiwSl3xW2PSChHcKzKxbfc3Dj96yT4to3urHspO6kJmu
jcBwZFxlwT3udj1LRCR+Ufa3Zs+FIjoW4R5KOZaMwmy3u4ZWTokDuXito8jgDjJgcN8bmvVV7bEw
URbE47GYqJWhXhF1oguRnyDaFL5/FfwvTJdnflQouPJ4kUrDfkADJhJfZt/5oLSlxUowCsWEZqsj
0vdq+HthXmwws/pVsrLD1OCWKlzJUP2SY/9RLTzN0Rl1Lb1v3CjmcCC/GZlSxBCq2gbcFaeoHskY
D8yplzCGk0RAuajkuQbQzS+EThgDnIVNyHKJjj9FhkwvDh9YrvLLUWWCWUw6Ynk+hHabhPyMPj8t
HaS9hs3XfHjPkwcoeWB0pLENyf7gmAoFzWwWDKQHtMdI5BxSqINTFYA7Sw0K/yGq+Jphu8r+IuZ8
Dh7AHFBgeV4FkcWboU65QrIMtHmRazRJUPPjUg7oqgx1er0sZdB55jOagP6Cac2ZOn9a2wv7wCkA
Nkf2tR5M8CVe1FdvDAXRZbG0W8eSaemAa2Bm7usZMHKnp1YryaBhVF1B5iPbjyqHhrdCwr5dmmAP
RsT7yCBbaPIcfcoVC9YRgQiV9d4v6TM0hvWkCf5zm833U1MWJSXHZ74VidcgmNThB7IwpssOs/7G
l+/KUSQiO4GmK6jfs8BK2TdUI9c3qs7z2rsrmqKr5AqM27+7e/Ab1kTvwUIQXvO9PI4TUMpNgO8u
A7GZWGIP5XdOZ2Uct4e4j25y662Wvt0hn+bcpWawhwLrZSrB0YdOAcAUiq1kvGKRc9/MowP9Zn4a
vZDLxzqpdAkoYf7AlimfI6O2eLPecOuoUO5UTtEyk5gXcGWtUhjF0p3ud0HUENctbgGoq8IgZhBz
1rWb/mPoQtU5r4fIDZzdg8zqZT36miCR2BzwWID3AjwyMBqwOqBqoLoTB42/YKc0mNi8blD2xzP2
VlDWUf9t8LCV7iTTHWmc7WztJGh4Uge7EU1mAyf/XtQJwZv+BB1ef5IS8fVLaSTQ+jnv5swTtpEf
U+vZMAw+2qz75c6iIbsdQ7Y4Mpbb7cvnjAE6goveOjYWZl02CW9Wvh0sWbfhuTy/s7JXrl5Gh+O3
MZyXzENJcA7JGhT3qGOtdige8bBDFKG/Hdg5lVzJGD0jJ9Z+8DXCq5vdSXkwQGOArkWTJM1bSTWB
zDaPoHMhI7j2rbqR/jPccaIEq9nOKMe6J+pkRs+1Uh1H9gIp4dhHhZbqVkl4qLOwmxDPjerUm5wT
Tcp+55HSqRt5BTjv1ajqFNbc+I3oBi9CiByCYh1d0i/SbSXeF4fPYs/KNqcWDfjlic4apSDXKF1h
Mal8/BBsQs1xcDCbSqvnVg+XQTRAlYaXcF1T0FSFak+WcaApmMCRU2q2B+qtYVnyNhq+33hrzRjL
pHTgCIGpVKOeJsH9Nf/7gb9O4Qw2hMA8jIGCda+KQIFJ853KWtWWkqFx1s+n1z76RWZOaR/fvaij
B/mMofsTScUVbwZdc6SI4ZwFG4YCYgWSsTdsltXjUnX+seYafSaOybRiUavYU6vCgFxNU7g+e4Da
uTM31om0G14kMc3Ts15fFxUpBo8l96Nbp5N0NnRs+jEINhCKGK5ntBDPAgeX9dH0GzYQM7hlTjdq
8j2cA6pJLdL4hdB/w5lir+wn4+tMXYGvxUOaayGhlmGeQX1pAr7bq+zsUkiKuVOJgYnlwBlNvjxN
aBGCl8sMbmUlBcEC+pMseka8YWvkduIeGfSCmf9SL+SywTaVTbKrFfXAccIJ+PRweX7csrhq2Igy
h8oQlyGCh+ojRmLeLMUYb3SBusvSiYuRNVQnppmvFRqCdc3NhbsZHZL5SeabFDo+wm9ctr1+iliP
7sgdLuA9et+cfz6Qff/QlC1EMBUWDMwECxnn1JOm3Iu9Izk0G4jFpcI9Lug9tOMl0LtY/qEoAbt6
PsyyzYMpraeLHT61URvFAQZSPJrox2f/H5wNGpInz+eADNK3zrU3TFols3wEoMwdUa4iV5BLAd73
KBUhxOa488fri+Op42mosdeD4xKHmf/9PB01IqGy7f+V8avaFNIQD9bhXsCWb1t+RYpGa8qnJ8O7
8W08cm8w3oMQh1rw2vRrZRfvaKyWCUTlJ1XSSEGgYjzPE9eg7t3i90xo48DEpj+nkYEfzIxvysMc
spTm7ioc1443M61D7pgMjxNyLhqqgENoZfjyeiHKZdJFNuHwt5NH75XmbgQYWalJ2bcmKNFrJuLG
ETa4J4Exg1j8f+1de1AEIopTzOGmNhIGr8fngrO0s6D6ohR5dvQMHzJgH1ZnKpEAvanTKab3pCqo
8LZFq0PMFgO2ruy28Lyla8FwDp3jsaTbv/qigdkDamnsZlkvd3St1u4wf7I2oCAlzW+yFOUxEXcD
ENLYj+rIlYcCtJUJZskoTPrE4rRX6gZIS8a+PLf/dL9UiAjoaEPB1Dypdq+xgTv6O5Gs3oA4nqPj
0hnidMiO8aodvf803DFVMDOBjIj6tlV5ZopevzrrZSqnWKpGXvNImNp3BFWlcANVn681wOSGbio9
wD4nBetb/bIc126lErnHohK7N8sxZltHoKGWBMW0IzSZmUdi3xWwOvv0BqUiNCfTlVY0qM6ipyrX
N7TqDLyek83gxkSq9ogc3LAZkCXoWPph++AdURtcyTm2UBebEL/Uw8m9QuqmddRbKxyoHe2SLodw
yZF5uot4LaGHTSCoCFDxb0i+rtLMDkVU7V+vLCBI4Bhd6wYhiajz/3oznPjp1Om/KnnarfCB30mz
/2LJHwFlYTrckJeHf/Hsgq6UUUBGF4g5umrQo4Z8oEzuvS7P6soGjMJBmbiLDw729RD7/vQwWJkF
4dYpIdv6ZPFWk8qI9UgncKbjzMV4kQtsEtSnIjWFWcZVZMZULVMayY/k5t4OenA4KotJ+Dsq7YBB
INUacP9Yy3v9zfvKjb8hDD6hgiqt1yzj6v1MRLS8fdePheioWUCuwuwbKYGNOZTfpBbkThg5IchK
kYh1ab1Z+JObogi9E/F0vn8SBwtUgfQys6LzbeuLJOvEtYHkQ967QIADYYoboSxHCOks22JSVKdQ
HdllVkE3AGeYdHsvgTh2wSW/1dljooUFGnNF/DqmmB8QmMQ02O2Srf1H136LqlgHf0ZFhix6OS9J
W/Fk4QtN2v/cEG3/CASmKFTUpXSX1/aSHbDAiL/U3Lres13GYlk2o5/C+zF9z9G2FJM7YpjJeKUB
rabwJ6zN5Vot5fj8r4KfFqZBV/UxMP++Xa2VlUPkGF1kM3TENQ2ae8A24b//wlue5skipxZZ6lQr
94mPw4nBKjP9xD7ULCS9K4cuuK5btMDc6s8H/Pytcgdpv09W+udtFrMKBr6uBoequy0jUUAb8F0Z
MwtCg56iM4vv0UepTE38+j6m3BRTaK6GxDW/CytDY6tBLWJKp+Af7XO8P8xNJCCrbiONyzF8yEC/
6EMcIbW/UGuIzgG4BKioVxRJQz8kUsmeaTDw7WxVhaZz1e98wQoYH+NePuItsHXpL7SZTXWFQdCc
xX8zwbtx7l2nvB4UhYXdTZqSgpza4ZAjaQZ3VRbxRnBXD4Wgr2TSJAaHkYo8tQBhCOjz8tQdCJKZ
9QTb47+R0NUg2MDvGHAvvTLV859D1XBnK5tuHGECt8+4pyCGBGnF+hGmiHkUkTWwvVBW1PHK+UWd
xbsjiggWh7961GXTotAQBePmiHFwp+fkA6NerIwxpYJpS+Zfjb1N+ZMVh7Il4ZvoNIHLIgvxPpPR
JpagNy8OAY94uMq/B18QdCtziB17KzkPfuYTz1ZeuyOwwhJDpNveOr6U548xZHqqG7CrnCW/zYtL
t6YcDW9Oc8Wp+JwxPlhYYvM922lZIErVr6slgZUmXHi+BMIEnFfw9h+ldG3ShgcANUjbbEmH+Xjt
hlsFwyH/TaDUv2YfnP2nOUouZJpbk3Mu38AqMv8iAcdj0UChWZvuhvFG6p/O3Xtmwm6+I8n/sfpW
OxnoJdI1isgUuNE4IwY2zsKE8CttqZ6hw8ZeOBvlDy1V23CkAmQpxUPoXUjAAZRceIoASOrIBCfB
1B+/8XbPu4IaP0TL60KxfLV0dNcgLS7lM1dn7uCUx0T2RPKSV0omqfBFJGAcT8BKUCYdMN/PyRQn
zM+WcknHQ7idJrYKiyI2o/er//TDEJRI+nnURJyTuLmnb8dspKIuf3cuMEik2gFjiAo1nAebBQyS
Ni7TEEfx8MALumyUxCTa6ly4nXRNg5ghd92ByaOCGUCKG72xPwxUp8KhA+//gHs19xHkOdfSdIpf
X+hBcSYxkeFYedYctajc7V/2VUs9/ymx49qjjUUPEertrYgmz699QVVpcad/z90Ll3EDRLvvpRFg
S2iAg5u+E8eX1Ijxz6gmKmpXvU4PEbyXklRpqEntBTmiRsFiM8vBAMkLwYVmDWzI5Ubmvkgl49oS
BhRfqwNq8wW+Phj/nZsc222DDGAuEyfpGW6jrd6avDH9Z1Sd7rUmKOqOW/XzwM/y4/7EpiRBRe2t
cKrYh6KPqlWKHWqPJdJhIOGJ2W6Tws23tbSjL+j+Yep7EEdKxPC6RuzhBZGElh4x6KqhRXgKTlOs
xfxg9ytNfnmGmG6ps+XmEvAlvIFuOoxiFMOolYQo9RIcn+0lvxe60NLk/b6iHWJiijR8WKquOiOQ
kMIG/g5bAc3v4fYF8JFeLvF5bkekK19isnQLEtYowC9DVi/fzABEkzw84T/nzJwr/ShJye2SxvSA
i1nmA8ZtHgGC1DrZfJxwGT1lsvy3ZRw408UnOhC87NTKhrPM0PKKXwROKZ1+NFdsopJwOTZYkcdX
O8nzWMjNEh7PXhS9D7hFkW6JYMk03oYprf6SaBmHNO6t9dqJpAzhKbF1inycSm3Y5zeyw/7P3c5n
CTC4F3HQNWNYjV4o/HVTNOmyPPI3DD6wRegqnaFh6z8HgUphO01D7NbeAV0hg7VSGSBGkfwQAw+q
zt6c0iORjsv/RmnlLEXuSPi9BbPtTQzCm+slOZy96LLAyU3MlrngF/Jpg39rka1JKlCVEvHK4jh2
0yPYxGZzcgvyPYNKG25upJ+1DQoVQEotaQ66v0ljAjMrLXIFloAuuvmUJBKSdcQQsqAuNyu1/1L1
eMZsyvTIFkn0ieXuniTgoHlPQzO93lRAbJIYCBfTgEUkmEBRk/NhqLU2O14miC+K9spLnYXRDjey
VdWo1fnGt3DHj1k1pe0TCmovwu3KnHFoZcfDN5r1PL9iFiSY9lFN1WCdcgCQXEBogwnXRObp0wIA
Oz0QBpHfOzyFCeTs3CY4FDkSXwFSAbQufXGYDdgOjOvC4EGVaY1yxEOYQlRH5TKNk3b5g7OuJPMW
OmpJKjAKCyTD3NHV2KvJbsTQMgejDH3pr/rKSMhGB50QLrj6wpyDMXtvop9Kc7feGIL6OlowQVx9
udlYFldD8DY08i35o1gl1Px8hLyHrAdNEMUjaA5STmhfKsWMtiDxG06I4P68woxaSf+oEBdasV4x
zr8ub+rL4nHxinF47/jNzWK95qCDv803bSchyv6OdK3U3g3/ykYpZBhCq2crGShhxmD70mLU4pFu
IOQ2K1BBPu/hcjRnU8pt8x0eQOyaD9dLKRwilcbyTXYu3ekS9konRQ7q5WaR9Ab/WMQsuc6rPxF9
C3HIPDmsx3QemeMKEfOzqtHGDwY56ceMG+3o0IgAWedVyadar7+I1T1h2JaIrP9fhloQhbMceUuO
3y4HWaq3X9OOnQQ549Br8R3iDY9TLor9FCU+nuKCO3xVpvSvgbaOkx9S0Br4gjcU2AYX0qcSCzzp
e+mtwZbBjySmrlLF7SGZRMME5PhT71IkIqtg4GVd+RjLQoFKqF9g3L/Ju8G+HfTXY2hs6TCeOcXq
IrwbXgFoUD2pWrYCeSnE+Fdv3+wGo2Wosfcr5mBAoB8oTaiZT0q3acLv1OU9Gk+X3zZ7tVu9piGf
xFBychE+VUl/vsNplWJuzGEdFWOubNE8MZd7c71DHKj9bKkKkmdtbGZhK4R2EF0i6126cazeuY7m
uzp1zzQlJkGeXMKqaoESlG2w0/hwtIYy3SVTggd7M5C1gtaWvHiJO+LizZ/EfkLtyAgzpqQ51i9U
kZjN39GnyUCaD96qLpI4b1JxXdT7PWrQNW5iOicU/eni5csEThaTE0NK2rSm/tWzoVUkjhswxWHW
I7IDUN7ZF8MYmeNVqb9qjUppRqPDrKhsWmzkc/6cLqIroMTDjceMyw7fa8pUx6HUwh+inLaTBsPi
pl3ivxgrwaSoF98FDJ7RjEDVysIBtNwWaPUTinuIZp06WqONbyZ2ix3zj0ZMqionTtSb4mkJ+Xa9
ycUnc9cPBymgaKYbfyGKYmco21jIxTo1SRcriZlJVw120bQjHme5hORroMjEXuNmEOY/K9LSzXry
giHUhCXEi8/notDRp9Vv5lsQcOpiAo8eFnyd6yMpBDGU5+nHAoToqk1rJlnkSbzxuM0sanUpoIyA
3V1TTovoH/b5kr09fxzP2AZCzi2qefia19oSw2gEJBUE67AvjJtr5UrwvN9pRSIBhwFwf1uj1DgL
JrVoRqaZ7dxGQ4Jl8FR0jm8XdVUS7TPiEXzMFxvLGAVBJ3LQTL2XPGAhO5OKYLvha4O71+wfjChn
GHSpTT3siUrJwd1ROokKBX1BTLYlMd4FV0oHoXTZWc1zT3Ei3RegOYQxb1stFwV57/SLuT35H7oc
fAw+CxsnU1DfE9ADSg8jkLufzj6QC6YYGGdKknsjZFjosG35gAPyvDYiAdrobyshOiHh20wNsR77
eUSb4+wa5WYmH0/YOJ/3BE+dESNop4SYP0/LCh5bppjMS8zFgkfpd61OnmHGVyGK3ZCXbV02/GMV
cX3PJXlr6vfcdW+baEuBMa2tXtC3pXoouGmcj96YEEgo8Br03YsJykSEV5h89OqXg8mhjUYc+/Np
7htADBurx5NIAXO0P8S2ZXlQ2iwlg7Q80F/sTHKns157NM5Oakq1Rq7jzzhPYNy0WNi42LAz68Rr
N5KhzRGXT5leWzJrdRNPL0LU5Rld/IfIZOBSApB9noyHzm3SYtYdi3py05M2D20PwMeRC37QWlZd
NMc8P977QvpV5BaF1dq0HjhXQfPX2/xVyjoATP1Zerr2MzjW4DDoasfMotSRE6l7moLgTd1BFOha
w/d9xvUQF+zI4EKQTIKbaWuoKS6YbpPMI8TuthFgEgNt2HKnwponBQSemJjFjehrq66lbrEzicrB
sH7I2AsFDOkZDIpo0KIuVm4wEILSIKrrk+Zp1xSicKU8QY/2SylDLZqiuZAAWhe6ganyOlEPFMFM
7xccxbmg0t2xRLSVXAsrfCeq61PHYyZGs3Ec/UDKEvP8wFjHzn7+NJCx9qDXcRQMy2iO/PSkGysl
T4za7+am56JQLqqVQUr3a4P8FCo3wBdAM21ud7JRdysDUby8Rdt7tIDKvo9X1fFp9YDPctDfp6G5
anHrq8f4t/AcK8+bxIMCmVFR6qSJ2V+N3BEeRJl8D2v8rp72YLikv/rVr0Yn6MM0ysrtkvs2wSMT
0WZnpmBvtjKI6cGDalG/0SYz714cMeQc4+D01UUGjFVBQAFohZ+akflx5Wx+8+abZrqVVqbfptBr
NUmkrAHeOVBp2CTN0B2cP5LlkQF2yBaxVWj66kzMSBeoqaBQVoV88q0N5+jcPFZhPXqa2RCvJKOY
00pio56s9+SX9xIBCmu/S5SAY2f5A9PFquypNYG/vDv8N/Ka+xYmqihkKTgabU80qq9wr7dJAW7D
dbNe53+MmdgfZlgJzxiAQiHl4mrIorA9wJRaijUzzYc3k0OPE0TsmTuoISmFLCPmda0R/w9jenv0
aRsQNWDGtx2ig7DbxZcTbI/sfxEFv51X9drafb2oO4e+yElrSlqePA+ZS3f8kgntTdn3UfYy/6BQ
1+Nc+ZZp9S4103PVCd6Lz6AKRWsgCx6tcKBK6/Bn48oslO/o6k/usL2kwHgOgHW8/vVO2lPFm/uw
XCchmnR/MfsZtHxIdqCRDLgcDVvDb8f2+cvte2tm+DGkcJIQRyajs4nQZcNSjWRa0kvUF6Bh8gbc
gaPbPpVGkN2B0mPh3u5ivg9ogH12rSItGQqySCIT/a00L/+ydRuSAqRfFd7Bu5g3vHLztR9kxtJC
EUBoOH2H7gKXs9D6h3AZNKMdsw54/zCeE7OCLZGGdh1861QhF8I+KeidE7MZgQcqHcy4EcQLfgOY
9hRu3xTRiQeXgRyQAtcXDSfAF8bx4OOYM4K5d80/8WHHobcEmiMxUsQjYJEhB6gL5HH4ENUzVE4o
24Szkxtpv87q2uzT78jbpuF1p4tLaWIwDjwDe3CUL77NYocZBreZi/wbzq4r+7n56i3tOvrEgk/h
dvo7cpNt9zJsTfBiVdYV8Aragx3uzl9LcGVXt5LP0+haBK6J6oM5npihswTDjh9k38YhURzztWDc
xn3yo9KGqHmMruoXXEFVw/kx2WJ8EvhVCxxForChENh4z5eViTso2lkmD2munOoHq4KX9GVgpzk1
qDRCB6mqUoltKE9zyd1N7f5eBVW/UG1AhBr75ewmn3zD/vWiICtlJY1exZC5wE67UNOJJQby67P7
W32bbc3GBM0FvMZzWKrnH/vcD1mfBNICl2pCeLkletv+20jRpRG40MAMZxRHIfPukEjIBSFOiJ4R
5qY3tNOgUZYvFm0sDCqxe5hpjo2qd27crlqH/DYvuiLOOuQFtVosY0nBy/KwIFKqp25ulrQ5Bm2v
GYk5rta6l8wrfqN1r/BTS2dLWCvLtRc6i2KNhkuICBqjVcXxMQexCP24/Mo4f9JA8A9/78BC3+UJ
4CSG/aBfXKpWew4A5UFPn+0r8LgG5FIbv8XM0HqiT8BZDZzs3Ds6ANjGPgfNQFCecR9dePJVPdmG
2hl6hbAnrGnKkN2ApfJzm9kS9wA2Y0GD+dvsE8fJPJR6VcE+cE/hxkvKMtopnqadRPoSJoG0oaEP
Z0lU5Z96YGKrs7AMnCLuERWTV7TfsikF7bDY2eg/PhMuoIlD6MJoMxwUaXM9TNuCDCP0TTPgWjIf
RtMTwDyblfEB+vclskC6rQKRKtFyzv//PdXp5KZjjJGIWuN0WqFMeNRFV+s7BPX6keNGYUY9zDJI
MJyD+f6h8XytfP+PUFkUH8VeW5sPlMuYpBM8WE+LGX13ZLoz6dvl+tTO+/eTAtKpG46VIkcyjL2Y
j8qsTH1k8UJ3YuUeM6ib0BG2lItnqvrfz6XX0eLlU4l4TC3Y7BkCxidsaBWLIUmAbKgYGNYbiqaQ
LDkSHVY/+cvgvukp0OnQUae0rPC1BUhNEtUuFD+9jScM/QFi7ErUyA+DZJrTI0om8PWd2Dvs0R4X
HHjWydOyKwp4x9XQADv0SwcU4JeBAeVx1jnG468P/yyZy/gRrqypm1yy0OCT+v1rWaDHECs1ACnm
xIqqjIc30SP+hN5xP8TKcNmmLxxuqfpcH5XTOzfxZRY8lwjQAlgCRT80WLeRrl6XSQM6cADVV0on
MTgmQ4EQOyCCaCLlwhnG3J+NHm2XfUGERXGl0cZ3XL6xksXSU515tgBiXfQfVEpaa+klBLdUipY1
mERkSpPfPsqlBtz2d+dNqsWKTulGeASIF1X1qbn/MZWX23iG5MTAbQt4mbQirGx4IKP8wRnqFiy5
3mZ4goOznnCudIpLE7xWasjqedvajMoYfs++TgVWiFgmS1wFM7KYzPVS/yhNpwHkX3mpO8JyBexQ
jE8b2VOHCoyfv+UmawOWE/1I2Ayn8/MkxjPqMdkwufpnGNNHPGdcA7eQeGqxar7Wk/FcrniwSjPq
Ft9mZdMc1BTrAIvfVX9yJvXorO1II0w4L4zbi3DFUpZd1aI9uA7eKCB6LRZa0oUEcH9gafFgr05x
d/lCr6NxSpvfjvsfJGMt6lwqtQ305dCp1ky84asBfm9GYjc2rLmi1xxH4HLYfbueP9QX8K/7Csuu
e3+be7UzXEq0tJmbZNhn3pWvjsb9iQlptjZkU212Xj4l3GeJ/OaTDkfFT3ScVcN+Gem82J5MnOOo
RP3oF9OPsTZL/7Wfn6EV0Op0Ed4oupGrAnUI5gQKmAXZnZkUXJ3V1MOcNgY+eJBdtw7EeASxIuXU
S5jo70VXKaXxJpmrr+5wmgWwa0dBwAgU8hxgIzgg/Qqbsfh7uN5QDuJPDWIGCeFDotChAoUNFsqc
N7J5Rgel+57TTjmq6ce5Pit1QxJjdyIIkSMEPsHfjhv3ZJr6hjn5wtH3DEsYBB8+s0GgMZ6yUyIt
q+qvPYYLHYYhzbTzoQzLAn9WtlY66qJWWnnXkRmIlaJBD2SUeBdT1zW2ZNlARWUk5mce83wrFxiv
aytDm98eGa+GZIOUvGU16J+ti1PRiG9MnREvxOoTdegvp807f0Njs7Fk2cATU7VMJ1dVg2CC5cYh
O2BCLTbkaQ6LPQ22gBtVoqOqO2fJSgBaUPIhoAR8rrmJWZFqR+ABBtDRC5MCNqPvsgjjeYwkRv8g
toH//VvxVBS7KIwVW8EOvS2lgH2xXkChVlpDycrduGlKR7E1zobRAWk+4OFBAgxerrR0OEjyh+EM
Kjh3Ogsv4M3SHa7iMOMDwCk0lXzx0eOyv7g/vZiIdCiqQ35T6HNtlyHjDNEHsFsxk7x6NL+baHRo
FJHLaLGP9JnxERvRTzblWm6YGSuTVLdYfqHYLJah/mkhMiCmzXjUWs8piRAY4NyhGDlvbbMXI50J
xMEz4CLpw/xX6Rn1c1gz7RV2X0HbUGgMCROUANiYdZes41k4wN/OAXWkZd3DKv39kquZg1j3cvL0
UueUQZ4H1r6jmwmRXtc0YxgjhUxYvZzsgpoN46yz12BB4igc7q/Ortla5elnmKqfbaQbwvL1IeIw
fN/Muab0Cf81PJLx7w4JbuIXUZTFOuB6U+5npavMiuh7b4/X7wtsCBTLrLrWtICRnjcaWE/mXgoW
Y2Ot4tN4yADat2ksXcJRX/yxKXPmy1bJBXjLPHYvQc7P2/UfXjHPGUwRAHVC4WW+yaoN0lFO2AvC
nWUJu6052kGhIKybBAhE2QT7T8+TV+y7cLoBz00o3KC3d0TeYeeC2ZJ5Piv7H7mHEU9v3ICOdqOT
hlK3npbMg85k3/U2z3zfCCQPuJwUCKAbneyFeWJuCXtSooJMur4mYVqY2UxS7hQ/HR9wdYdLWOZn
1/LwSXOAWLzEpj3Q95FJpGLN48M996JfPsd/h7B9A7Q6TBtELcQGZZajqFIM2IDe1OKuO//66wN/
Fdqjw6EZoBXxr6dBUgPBA8tcfSqDAUdOBNbl7jMR7hNwXL9dNGOpnitsICxqOhLDhoh/nH00Xpx6
0qBiGkkiEvu+7Ail8Bl9S1fUXJ21+r5ARaOGOJM/7Lw3Fcv+KKHkdWHaec/gGlki8AYXNld3xp4x
PbRsQYsezt/tWyYtuKZeJavM90Vsm0xgjBZkOJDRGdFW4A3CoZ4BcxYNOFimNT0ASxJtVKQj6vor
yfjogY+sc46PYHgY6eaDcPb+6jTlUH/lMxEYVMylZzdOhsDEQ32/Gu8hQvWA9lUHJ94U9u21ibav
fACK98N1NY0+O8NNKyYPz/VL5nh6MCRk4ke9iAAIG3LnXm3x0ZEOnhHo5byDwkosNnQOu2+bMVnj
5yGhkfuW0C+54MhwMppRd4XYLM9WhnsfeFty8UPWmsYDOP4RUPzbQWoLelHcSVmEbnY8dye7PxFG
tiE/sM3SMLWQNdgtTckWuygzbjrZa1im0m8370oTTGE9e22ozr2G0z0+wQMLxuQcGSSKNt409FKG
/BWtdjOQsHMon2kOB9BKhI1al4DF+QbAH0Zsqy/+dPzVYo61X0DjjqrG4RHR6fTryWnmqzgWoeRY
Y+O1BxEY5fUETdKA3EN8MdBEEve9Kk2zBYX+yy9Kt9EstPFoxQaNm/hKMcfswuWVOo3m7bC2a4M9
QMhI4hrVhWpVhYTF75eWeymAKOiikhEKRoaptoinC6LFUVxglBugJN1C74dyE3HQy+nuMz7UJbL7
VzRwgk3x9EQyp9UyU2KWNGFr03frXkZKvIiG/poWTBy0IXE93j/v405unP83ufFKpVf8uBRsWPHD
eh9hW8qKd1ilAFUg0TlljeajtywS6MKx16wSIrjD/9Nkq8BopSkMcWB4u1RxWvjdb85n/mJy08ES
mKnYXbZEkoMU/aii953c6OiXMHCsrE+u9Uv7UEQb2f/I6FNfJZ7GPSroJBri4Rt0tuUC1rl3qS+j
x6m5WPvL58dtoKRDWT9bSS1aFwZXdOqGq6tqh2rC9FJgn1Z4Ur83qSi/9iXnClzMKz56pfJnRk3w
vqSMGrjId6e8BB5wj25SbulQ/Bi89XFb/XHLPXdGDnRm3nS+Crd4l3Sn/af1jaWFdzXgJiJEFSo+
jCi7Sln/1+nPtggJMiJgoBoks51AiKukqeHcd/zLMrrFncS2sQSIdryaAmj9v/5v0Gt7vvSoPi0V
OEMh3m4te7sYZsRAO+g920IJYlVmSyRS+qgmLpHQZwIx1QWvP7kJPfkDhdSriKEDG781fyxKdKpS
dFmENRxgy2Ie1RIofdNfntFfmjdP02/dMqtZjuo7cw+Ogk6JDXSuIJSQAyb2w2wRBYF52ntBz4fF
wQGBDcC84Hzem+baPz1vS3mFizVRK122/aAhTX56Wmpn83uvcxhieINJ7Z/IeWICkUrSVZGqsBJH
SXehMYPXDMYTd5ynIpqIZm+QX1qo1TtUmuCR948soRXaTvaS6B8bs2xfawu9fIgk3C/PhBXnWgtw
3sO4gdElRwK86mwq9Q5J1p1cZKurLIqlSQ5Uka+z2SpTvM4YCqWpLu7KbaN4B/6tn9MmL9D8q2o9
Gl0GmAxsm6Uhv80c2VMLfBbjBhGRM78I8Rlt7JhF3J3pJyWVHJrga4QOozFJx5LDcbx7LZtr0XHH
ppTnQHrmO56dfVxXNEC9PtifpB3YoLloe4A013wAsLkfa6rfuCckmtuRN1IAejJSZkC6+qvWcXQz
h2Zs6HfHd9nG/K2V++B0vSqy8j9c+qYfc0wwKy3qF5wtUWOBRn8EfOp6gaZwbAfYFLPtFYGozBP6
KLW8zz7DUhtNmL3ojtnaBv8MkYJ6JST3i75YEj+cb8ok9MNMMS8bWhGpSZ5lq7QKZzEgaHXjn6Ot
IyuFRzZT+SNFM68UapGdimyQL+XigPacGsJazF8GdBvGOxcpFnMXQcVMrNFcC5SyyAQvulUQmstA
2vtuGZUOVoPjYRMVEMNOY9cFs6uwzohIjD2WcaPg69ZWrTupf3wsa64QQVfuE4ORlae1xN88oH7p
yIGhNUcQymYnWfeBvdMthG7kd1aUhIqRc/Wt1Tdq8mxPIsCynW8GGpLygd6BEcZfvENPni6XIsAE
5QTycubTvJC1iXOJZ9N68K2byEmG2wue29sizXf7fYRoZeXTfjEWXt3igSsUQ1ruN+11smCYmkWK
Wur9VT2h/YIezuOED4tTrtdHl1rx36PC2dDScaXZkZd8DZ64w4VMxCEt5I1mJvb+MU+05T+VkfwX
NhAB8pawEBhMzmADrZQi2KE7hIjpid6bN7S9SPOQMJFA8/iaC+54xIflEioIfmhzwQ+C3fMYvKUW
LMWqL0UW9fkxdrNgzHHCIH2l+4CXCzmDtS5B1wHqLq7s8Tsl2TZJX8+YT0JcZ83XtojcK7hRAocO
8gV7BnjkLb5QubrnyS9q78ds5NLnNAB2v/0ZLwyUThgjSW9FW8a+VZBHG588swjno8G4VPxfYQm/
+2wE/JbDmJNneWSJMIhNoqhk2z0UJCM8M3uYMGxnnMM9h5RVsgHSMqftWgVSAaMNxkvJUU8iM3XZ
Hy68RXGohaz6DOx76DKYFLeBjdwja0k6n+PAhdTtziPHtsyjVg+NiZnmCGAwNeujlbrmdPA5VJJ+
o4Ju3g8W6b/9qxestV/sYEFcZc9kpOsWg9AEyq8J8QSGnjjQlmtzxEke/xP7Y3qGpas/MSMKZQK+
tGehMyAotgF2op2LwNA5n9RMBcJWRZQEt1C6irtHFRayCvxG0K2mDgRZ2YuB0JdcPtt3p2C2X0Vp
5eLUI6edRyALFRY6e84jjuB5Hb24EtsEIkciC7CoIDbcpuPwUBVvSoPj5gDurDMinwzSVYjFED3V
GH1VnNUNwW2dZQYPqk8qczbo+wmwM+o+6cooeCCuS7XT6/lqPSSY9slgA9bk7VGbnpNvF3y2IXsi
uEc9gj/e/v7h667hWkVWFV25yR8fGI6dBO4Rm37lYBsCXJy6B9P9APi0objXTVRkrGeKJAmAQlVe
7fiIVtt5UZx1olNY1oqyx81xrx8hL+tuvhCzZLe0lL5xpWqLc/MD/Tm5wrmUuTFqs9j51wLzp/3X
0/4GqmaaA24Q/Dnpt12CBimxxeBkNVKIbmIOtR2nuPsEZv63S2BfQ7jDxAFcx/GwWzegE3xMKw3Z
XuTnsRd6gmtshlapvmmSAOjvc6k8oMqpHoSCan0QQ/X2WJQTawAm+jTr7gEJjxjIvVH/K+T8I4bv
5s+Qrn0TlFKj50L0RD7buqKQ2jMMioSq+Qevsl4w9idVDl/y1nyktSDAftL8nyisLX6F87O3R86a
BqjHxZC8Rst1K0agnpt2KjW3iRThoO90xKcNv0gE+LfYyHRUwwXkDWfbFlIcJxVBW9vrEAAcaeO5
xXoj8z1RwyIO0HueZYjgVgDxRkyZrYiEEnXqm4OjYjcPEKugdmXd/U2SH2w3dpoMaCsMphR85OtX
/yol3j3/tG0QzJ/Qm29LaR75iM5osmmU3EPW9aIaVFjDu6bSDoXakeIV6sXmyYAAw5odWDePISA6
iyJCClihWZY65zobVdd4w4PuBYiOy+EZspPGM2cR+VZKmF8N2jGoMtBpYM8O49zOGscJoeYDBQ8I
PlMK4itZHadZ+pmOL9SyetL5pq+Bf7loNLkZ1MP4m7Q1UB//FCZmx8xWmrVKrU9RuxgnLqqiYf/V
mqrGxiSdDEMtfDK0eOgdEWFHKVRS+EqOp4zlSW1uK+zWMBY57HT9p2G9YLClQ1qZi6ECOiVzPAkd
EhiBxVphNK1OabknyrlJOwxOMq07TKQMU+AzuYSATQKQ+xsCcqfNvNka1Jf98Tq43/CSAK/AvT41
VUJPshEbUQCu7bd/zx5qODhyncXp159D3PUpayqC21agGNEsiDYSHSP/25zH1V+FChNRl4dQEVxC
24U8AWnjqR4tf1qBQGkLFov68OsZnij6LPEcyP6BL35wgax685yJdhOSmiLJ5zzrVPa7CyJyWS7N
LhberCTbiEocZm6CWlbE5mEhtjdymPkq/8ZoSv9++XHjAtHSB9bQjIWwMNJv2WO9N8CwPmyP/ach
c7HW2+FHwlQ2oUIS5VdMSw+ywycP40Hyj930jIuxrmHFe2FZJu5+ck3DptSK3Nx6RR5RYSgm7wLC
o9hJ+uDLAn8eFX27X8MFcOl4s5llol2yLN7MtjmVTpWtPIkuTwqFvjXWiYhL3V6DvB4pzWoea2NM
SpU1m+1bl8PXa3zOwX2iC742vANByXVNIlLR4QZ/T9G+92HXFisa719WvXOB+a7yjM5qPZVTvPPS
A9jII/mdu/DdC4YfP90/WLoZu+cLwi5cHQ1xCx13+Xptf1+7487DMJClHs48sCVPb8jDkv/xeGIf
sLXDIm2w4W1Qc7J0EZjrzGWgkHMHELRXCKnQzCm4HNasGJnlRFns1ZlQYb7zcIqLfmqrCehRI8jK
0gADiTu+RytwQRK3dYtFxZX4zuJOFxm3nk0ZfJvXH843OskG6z3/Lk+awUOC726lD+NiQNL7zewc
KbQt8wtBX1ZMPqEA1743Y9hXZwt7LHa1fZPDSU+e1TQJ8H5eNXaTpktABUFcCTY8jrP4y2G/vmQ1
NSbtqw1kLMUkdCffpr0mTZCxnQTKjQSWYvoSdjHz+DHYPtD7OR6t3B5pamrLnbdq7BlcDGUbiXzH
dfcQ9birc36+qXdqe3+KoqElxKJWzYzMCw/AeSiQesFnFCNoS4+0GndmobR4tYMJWqdMaQw8b5Lm
5hqEXlo0aki324z3vBIAYQmn6lFH57aC+6Awp/YmnOhdoK+eqIMy5YPnmmzBVDfWDdiI/Rv9kgsa
MNT2fY8THEm7V108MEMw5V41UNWVd0uKqCdfu8Qpm1+5iGCI7ywvbHPunlUQHe5Y0fP31Z5qpZ4k
AWDggqR8rqTjDDO1PsONSAIZ8oSM2it7vSLja2cgMrsWZ+KeV0VReXRe+FlrKG35b8Hh4H9pS/3t
Awz9ae4ITJceA5TjNgHocikZ74zh6B0USWU9B7gDg2mTRxEKCaUth4YVp/LMJvw5HX1b0sbPJU9Y
Zz8ZLmUnVxfl4F5eahJXFBtQtKiAOcJycxE4BSoswTonqouQpb6jPLx6quEpV50hbgGuCuZagB5c
j9SF5IoFRpuYGvGVu7fHxzGIsvPvtgSCR2OGEAICpY+hMIEKyykMkaFBatyIrrIODFva/mSy2amG
hZ7NFXjdrNOzSRnl89hJ5lUFjEvejyaDwcNYdeBcNS3SJD7IxHiP+CBSVENbqkCouwoYoYyzmz9C
6JrVQD2u5hWWGw+5kMTC/D5EcLxgKyckkrrFtzukgp+8sRiQtzxmY7ffroBl/0/dO051C8QeC598
BL8o4jZ3o6njhRTDwOqS6wJI76x+OhiVaE65F9ympVujXvHKYBXX7cpkIxWnRS/iIIo4vIXBT0zm
XtWdCOKseulACad0yBGhYz4SJKziG+mYKmqok64Q5sYhNck0CdwKLITVkrXMN20wtI6s7wl5lxU5
xuRg2vGKYDZWri9Jjj4KUN0tSkHmlEA23535iGCcVCgdoDJVYI4zRVRvr/Av77udarGFByHeYGRX
DIocHN3VzmsELd6NnwTZEAx5nDhHVT4mdMj6Nhm6Qj1/ptF1u/gFyRq0ulRb1A/HI2c8CCmOkfEG
uBQUocdmQ34VS0N2jx0tsZQ+Z8XexSUm0HJLhHlFplThqgBR2Fp8aabxLOnCc8TxmaFIoL4iSyWQ
SL5gSbZavT6Ezd1H3QmKM2ctUK2BMYgjwtC3jZBL6GtUWvkWQeIoVMFwCIqJbBZ9DcWheHtrH/JQ
HG2qjIVQZjPCVy2NplykJbfWoCuk/mRJICncbgfH6tDZ61vV5tKNUVRj6iLoTYywN81XYTHmrFeq
+HnWnhUlmGR6DERzI7/uMzJujVfAxC31v4BBnF38+wJbppZxGmjLAWmlg/siQz6KbIxYOo5z6yqF
ju10qjitXEz+qeU2rmOWt56kVIstpaLHn1EEprcdKD1NoGrNZfF/RyFJsWI0E5/4ZmY6s+6EH08I
TX4mEMxGw07VjSuyoaRwTYfiZJggj/I6KypMDIv0psE5AdZXb5WUWplNmnoDPvcEo94GIDqaGPN4
0JTJP+w9S9iqK3FsUcYtt9H8MKY/CO8szbYyVWNFC6X+WeMYYhRgPLxYH5+zNmfDZle6WEFQWrfM
qzQtfnD9AjbmNxbimXroyWUMvQjIgpjM/jSyv3eMM/pnTARRhFKGves3Nqmxf6yzkCs4ro2CpzsX
kZuevF917YzwctK6Ck1ZMSp4Pi41OUiryfOWt+LL0A3Ujt4iqWXiPxwW5ZFcCSb/XiReafEF98BZ
jP5jWIZNWNdRWeTktF/rAQGTvttzTflGvEoecQtBYCQkkqBfDUdrm2hM1kN9mUEheV8UgP1Dxvh+
xBt0FcjShHTB2VzTvyOSmW6DrnDwy4jK9P7vX+zN0SZaPFmT7y0SUMJ5ERsvLVifGfssrC9N+BzK
bZlbRyRaA3ktTu2F3pJPVEeXAkwgtCjoPZ4q+XrYs+pTj+X3WVTfwB8KweOUJcUUiKF2QsPIYm3H
j4flqCaK0rEM4U8kP8pW2rrfIanEujTLBsVyF4nac9HLMt29ant5aMp2hmMtX7iOqZS/5P1FN43Q
5kpNCXnRkYhYaS5K2sOpRpskJ0YAtYhrNM3t3hWaHCphVBnigPr9OUlK5cpAgvkHgD9RKTAxWNg5
tMbIjLZJ21rxV0AL4sE7x3VhZDqats/spxO1Y2ER3Bn9ZisKlB9SxmBsSTBmTO36rMossCPI61fe
hvL4FKPmAMf6eKlzzoCU+wStKkQ3f1+8y+71G5lNOBAYlgU8sQLb/o1ri0qkIONxQLRwIewLIekh
SW1ffKZo66I1Mb4gkc1g9tgo8+s7d243g9eJOwTugkE4F+sp3wdYajM9DY5tT0Q9367rcRgI0W+v
4XOcySgJlrS5kt/PRuVSPL8xZHxs6PnG/6nZPZX24XofDq/aXuC1N58J/yTj3WuKKryw9MBHT2NT
WQ8vVsPb9UHJvrDF9I/8dn+P1TV/ky1eTKCYcij7IB3HxKFGjPXG5fYozXX7Zku8uiQggy2Erlnb
ApshGoeALE/LoI39f9syMDuwma4VWnza3vUeRCTMS9AL281Fx2vZfHnDLJvTmwAlP9TnpjomEbLv
V9ewC1O4P9RSFxXGsLCu0C7NVeUC2fbW1uGgd7bxZrU/spRDDiRjRRxMK037O2jw8yM/GC4R8d2Z
6jZAVqmYVgM0iMfrNZqd1m3hais7ny8IEr3S6wHBc0vF3bf7rmOzkoOXs8OGx7rS7yHVlvj7//va
LR2/RE1vPdPF+WNnBX9mHw+l9Hod20JRduKH/62mECpqGep2FW4sLeOara3LEhn0ujp3ti8Po2OA
8o2tqGiW+IPET3/gsodPBbzY+B4ZCOKuMhRAuC2zQIDx3t05qpwaB7Z6jEsyBy3hheCchFxnMRr2
vW30zN/aob9Q4N74JNfrJB8HTAjk6f6NjW0wlbxl/B5uzxcpBtqtBKywWSeooda+A4+cVvKaHCVP
MkZZSJfe5xe+VmY1GPsO7ofsM+MoiH2rU/HxkKuhdeHCVBm0OAj58AUsEMWnYXP/0S5fE937HEtc
XPM8VrfqAsiHHbxUhy3p+4MYUKN+5RoAKF0HNBWPaIfpHQrP5jwHhkCCxG6ucenF8V8T7snoAumh
Mf7sR5AZhf+Me4j4y5llJjhK6/SEF2Oz4x/17eQ0izW5udUnXBMSUrt1udvMl8bg0xY2cNmeoN+d
InekzvnR7UAF7JgWpHypWTnSu5GNNmAswKjUT6y2owjnq7V9hv7CXZRzXQ2TDoUqb8k6JsMTy79V
0aXehazH7icpHDVi8r08TYvBLo/A/5LAq/SJuWDPx42LPKy8S/9FxILaVd4+dYIvC/q+H7Kfukq5
WDPGBw5/J2YR0Bd44WLPjGRD7ajuVmZLvIjTyLsyKmcQsNymsAtHoiOXt54NjYh1ifjPdWywwUrI
+4kKLxLEdCA2tuCI8bElqz9ND2Ylb+rsYL9yJD7NCs6i7S4/Bc9WAdAqTFP/fmg7Q6626nern8Jv
oxcQtZOhwiui6B1nTn9fGoXQY9qAhwaSvoCU8h3Ksfwo0C84R4+1RAywkkMtFUNU/dfCoheA9P+8
/xIZRRRJ82XHsbeVGdWHeAt7b2iohigO0KQKt9CMoOnVu9xEw7yJKkWKCIu4d+RpcdxgD/tVHVOc
RNcIUeS9zsX64wiBaQ1huPbcgz6z32k+D9OHT475o5E5+Yyj9DY0fFpFHd4PMW1Bz6qJBGxiy1eP
OfPG7c30gXRC6JM5UWg06nmS/3SBoda7RJXW1OxG19OJ8rRg+ehOnkth2AHTnvdioyZxDMf9fWpm
QEnoTPT7liZOww3Gqz/aZbH8h6JJWm1layDh5fYnlCJHbEiTY23E9MbVINS35OkkfZc0AeuMYsLZ
cCQLk51ZQgbGae6m2nUtTSp14j6PBEtxqsRoj7DEJL4GujcA3q4fA2FCtTWy+AfGZI/Ot77c0tea
CNDcenbPMzD/k6W9ft2wwc+dbD4BrTG277CruT3hJDq7FxN0fAH+VDG/loZaNmYexTNYxnIy1uYK
PaMoW1xJFdCJYH/2eZd7r7PBfighr4kJa2jVeNd49Z+r5+Y7ghGwVehZykHZPsE1en9N9znq9seB
h0bWPqIRUNXgojmyoKwEYc41fdPVLT1ElCcm7j8cw1PACDx4OGTtLGQmKhSOcp0UWBu4dp3/Zhz9
ouZ9/pDN2mhCexicCrMT325E2Ny7mM8TsK2YbvEsRVcoMQ3KEssD/j4Qazs+Ws+o21zeo5b+Y6Ne
QbbXKPV5Gjv0tKhhn8ah1uABpdduzHsHMWnXyRSThIjfJH2YCCEO3qaM0XNVATdT5QxT4dqO+T8C
r7hzrlCI4rWTo0gQyME/sZDxtsy6x4aDJXNx2wKzgL/hjmYR0R+PJU7ZrS0YkvE8JYp9gh/kdKOm
He8uSut1otouSdjo733u7t1eVZz77+McHU9Z3rBJgDRdO2yFncCKfI3/OUQOtO4bTpk7mERBHP8j
DOLzaL9xA0LTVMwWWSVDJWFcK91k8HqqaDGjGdwnOTgC5lNvK7XHUGL9JEiz4h3KLAcvC4tMY/7W
iD0WOeBRZzs6a04LTc02hX/3bFcE0GfQAVxT+dMRJ53ELQBwCLogkI+5+2jTBKxD4Q1/Elbs6quj
8QgJaSl+FMUojc8o71gQAyd72zqwk20rt380PqLnhjE/3D790yP2f9jCjyO8tvmEY9dl+FNUzw6J
FeYUWDRrl6GEu7t48zzF5rCpUneMzXJ7ItHGjYlPYpcZWbEiQrqEBUvyYR1WCxn83NMqbqmryYjO
cIHM9IOQs6YxbQF13LgOR4H1zwMI0u22D7DnhPsBWWqULAHNo+TuWUQthKUsQAEM8rT5y9npXpBe
0G4ZUjaGwoRiXt+SUlr84nIW48eLXb/NphYd/D/z/PsWtzmQ4s+M7LcvHdEzYLGf1G/9MRtEEdFL
NlWyvs0qoKQuaMgl2Mk9TC03cgPInQN/EWhjCBj8I/AVH+s+sDWiFEWIaiBY0fythAvIDmX196Sf
lQJJ/HXKaNLrpgNmSrkUNDgQevoZ25ES710HQtcBThsaQYmcFXosg/eCzX8jMzaR0ngljn5Tq6Z4
GISrbpwkBtcRToW0KP6VOeTHMpoYku09YeXqkpr5cebXNZL5LSI8e9dslLGPKbEnaJj2crEGXAFa
YEIBzbrM5qQRPllC0NBdmeU/Tfs8ialhRnp+elM/8+bxdj+o1GvGCXtbOVZIDviks7orkt7v3jcr
GYVV3bAeoCv7bS//VCKawIkDpUZg5Xp/Wci6bD13YU+gaJiF6xywOxq5WycMU0OZA05H0XxxxgGr
CZfNV9X+jfhZV18Dxi1WxGZUaFq/1RZB2a3Tfs3r1v+SMWDsWtQlJmnQ6N593r0t+uh3GJBORnJw
lUZ1l4hapfyGtVQhAY0Q7vAzqOuCz25NNE0Oy2JThi7A1IeZK4RXbedyEKB6tnlCOBPd2dIq/2+h
woQXigQyl91gbr3ZFL22Oeit1ycQ9mv8WsLAEkDyHS7pmUOEXUll48+rhkLUTJrPDSbqlUjFByTn
dEFZkZP467WzDbpM7PF02YKFL9eS0ojC+qnNRebbQ+U5QtlMY51zTSlCvlMEPxS/0E/MJjCpEr6o
o4fB8Yn7T+mLv6sWN860l0o7sETTIzwI09heqhFfRfmbjGeU1Ruqy7oN2LsYfAc75i7aSEmqusA/
X04SwS9J3VPy9KWlwzxnCFfsC1BbH3LnrcJaqgL6hf7ObE2Hc8K2+SG9heGOo2xKQDEhHHBJRqFt
y13Awy821TEVcpRZk/UO5rnEp0+dY/SyBl86FnHpnlnWW5yuAbNGJS51Z6ZGntvNMBcoHPegDJ5u
ZjdjuJywTVq3QSQxm9v2A+zjZTl1dU0GEgb+mzgxjyh2ARvzBweBl1j10vKpz1OJ0clGoI+RGvzP
BTG3YuA58Ivj/gckitCkveSxb1jXrS9xxeU8aw3xZn5D+nlokYvDFrpik8/L/M2Yz2J15bdQUudR
LnEhjx1bFeEKb+YkFC5t5AF415zsecAiQkyG1mMAZ3Gi+//rIRf2OLKYxTqIR1A6UxYyp1e0+1eh
QDgcb+5VNH0aKav4UqLwblY0ZofOjNBKAHWTLZwZo5YODTMpGZ6KPCHg4ZvD/NSK0XnkGDhytgue
mmYgGji5CN7XF25xrLMKKdvBj2c4/Y39WaQYr3X7lSNvg5HVPvM00pMjmkJ2acxSWmGrWAYUwXQm
llFUltT/GGAQChv3M8fnNBCYGUXrEKL94RHt4PIR1Xv0CwzIdDU+DiTr45BLJzSafupBkxO1XLnZ
T9rurBjF76YjQU+YPv+mbjSE4S3YoNIfGYCgj0UAJA/l2D4qB4ysCozt2mV+WiH76EyV/m/u3qIm
+nEX+I6FDflR/WyLx7k0Grz8OrICdXeRH5Mk34Lx+098uudzBRmHLoECzewR+o45pHOtmbirHVjH
gJhsnwnlFTu/0/9IwNL6gFMedDJwUr6a5iugJoKOUh+fkYER5bg6THGfg1kixQy3qDVPMg51M2Gq
Ltz8Kp3Dvel1FnpEWiBQ8DBhihzXsM//ekBTcOudEwMVOTLDRZqmDB/BweC117zddVRaTlBfGfuL
LIYb4Gb3IEsjbm8hxshNE0+lcAkDirIih3s3mQnTiDuXZfEpwg8aXaux0BV/uDl481feUA7MxnlU
ZJ0fMGuKWz2B2G2iCnUGImvB46af6inLBNEa1bYP7XzMlbSkd0LwxhVfnSYOD/nC+jZ1KzYEge38
FLFaw+/SzK1XSL+nRhzkfcDLQwgnu6jGDdQhOwh6Yof4rTgdXR8Ezu7Dh6iuLdnESPlLOKUBBIxl
Bbd6XUm4fBFXcFI7nRp4qga1WboBQGnG7E6cxDNov+lkIHFZRor4ElnqVtesUmTgYKKGYU7lSLMu
U47vRLq33irvmAoi7oTQcall89Hrt4E05DOAXb72M8/7hjZ9BhNLmt0Ok7C2ZmZyPKhooBiZpBWt
q0WRqih+rc0cAuFH4lmFNUpk8ywwB+IfyFVz7AYU4dMp2a58d81I/fGeGgIP3gWH/nwgkf3ZbP1B
RN0HyQknUWbaI3Qz3ZTF/5bQ11Crfpwhhl/o5azwAjW20qWU3YUpRWH7OuIv52+pPuvosiYa3jJY
UthNGpJ4+ffB4f30wT+SiNLFvu5eyzJ4CKNSFxz6SESPY1hFky5WmcXjvtcbpv7alaIb9BJuPQ8Q
TdZ5+hOUvnvI4iywztWiFep9Udg+HGIulfs+p1v0sXWgtr69xnhbrMcDDT7rnzhRH7xIU2YZ11Cp
pccz5z7se77mSANZNoFPLlBkpgmVy7JJHQsIVqnzQ2r3SkIDx/213I4D2cfdUidK/+qdKXAtzRVL
qWdq8XK3MlTycUaxKlZjxIO/c0VRQy7PIoFkhKM53B9/TVfkcqmyP1Dmb8J7FrT1i1FZQ8TSYKbT
kKmwCjTVGPaBTOUHsBgZPXwcZIEeQvzlFBx4xDxaUrJubLDtoDkTHeBhzpJDEL6/WV+IAeykudEt
fa3nRJls1O4jDT0UFy5YqiQUV+zTK6ybQyHZ+KMmDi7fxmsWfq+saCfn8wsd2iybke7H7i4/I2CW
m5fpVtiUFQcjXIAxHPvvKqWp/DF0R+BOQ1lMNvtX7jX+m9hYb8j5IYMU68gy+QxhPf6yAeQAa/yu
hSarJBwfVPJo56bhZbodvuBTsSgIOo8BbZ9xZAulkMeEw4kRobipAUy5QGSVvaH9ECf0Y1u31quW
Zd+Eaz6DZQdICXBOoGk/oxr8UWjMgA1ACaFAcedR2yO7TVEX/QVijsI++uOV6xl+tWcEKISN7YUT
DZ/nsbHk7APSo24hfac1eA7yLddQXD4YtzRd2gnuMh5Q79o4ai569PX8ShwgaQIaMZp3bEq0Ghkx
lTmnMOZGRYk/LsQGnlSIjz60jfdESffsD9in1ZiNSMf2U2CSoCfodAnsVtkWj4hiUEw/LLWafU6f
MmCbRkHC5ajMibeStIZ6PhKUFdSV+BtMNM1tt1vxLJX2xJn5v8LP36EXpaRmXocVeTEbWvY1flf5
YJCDctYe5rYhLeOlN63IEFVBVlH73xpD0Z50QuSlcpAY369znv8Yh0MkLhlkQyzhEHlWXsSkGwgK
C2nFZfNZq9EPuFxBSHxAFAxSXwKwJmkghuEA87NEfmLEuewvNlTqArhT1D6XqzZpFTklSsMm3xcb
tlDohwgDgYdOlCfe5ufn7WbDlSixMJzK31RtCzooWrwnvZcfa5shBIe+WuWWNNwGJPzLV5u/OjXc
3YRlBBLatKrQt5nCAnDYeldNnDR1o1+qMzukrNtlYUSSZOI5bFu2lMVYLWrYD/2g3u856fg37ZWa
IKIK5S84eV+5MclTHsc2PbMvQ9DOd35MrBKd6GZkG0KWG+TV1P9wMGY+0XYqaUgibpvtelTX91Ph
AfViqpErfmpY+XjPSLUtJlD+DcyFQsOdauJAlS4eB9e2+JNuxfbFMS520WT5nVHu4pgmbn/V9zHe
mLcLa2kqwCKVrg3G/1WxLwbZz51txBVQeBO892rla0OiAiZ/DtIRv5GJzB6VQhlc4Wj8cReXnq0w
NGB6359Ex/yCnkwzWOWc+cgePxrtqedLMMS9X5DgINf8z65JieUpKDq1Ubi1CGwDMZ/O+UbGCki1
yPliD7Jgu+XrhWxvlchjjLVKvci8GAN+ExoUHLKCaEN84EqC4UGQZbccrR38u7Udws7f7TSL0id5
EoiZxFo7WUttoxx6kcgIsg5C1ddlD12IVAD3JroGPgUi7cTbHUL3Ruxj77boZLMUDfuhDGp6SKsV
1KXvi08rXtW0Y5zmVs8H4Trqet9RQXp/LWVY4GoVRUhypdwo4pOy7mYCl2qJ2PJEc00/d3GNskER
Kt2Kq2L9K1jVIpC66l+kZbpPMrfE/zN7ci22wtZ2YIB20f/LR0zvuBM2n9h9YI5DHO7fdIP9ZOuR
SyTcaCUzTw7rvSHFrWUG68dYOHhQdoXJ4GcZL8QNLJZBfIZuxPBiDrKX0SNlOlSXw8PvZhdMlMny
VXh9kxgKsgpTcQc9+vSbd9jrTanA3XVqKxu5EM8SrtuhWtuJOHH5Y+pduVZ9PB2mYyfVmD/SS5jC
YL/52G5TcvQPxQI+z/7lIW7ieCYBU5upcarKZkE0jS/qBi/HQgAIF5yNS1rw46Au5FIM/iJLDlB/
MJOvh5WNDm/ucUL07H7MWwI9vCbA+IrPtW4/cLPZMNNUIsrVcOANQ9dYUMKdkNgA/H45j82+ppsd
DpXfYH6Pmc56iDzpzgQOXVxIf2p4vV2v/hqGt6xuN9dVL4VN4+fqW5WnUz9l0m1e0xJ7ZUAB6BC9
7cQiXbFpjxMmKuelSdMiWoL4wYFw8BPKMXtzWlj9y05yMIDfE8uU/ExPgVqWIV+/3AfZIthUzxu4
Hj8/HyMMQ5weAg49SUxdVhWqxghmIb860DBoQ4qglvrYokz+ADFGRKasyjqtyrGY8KGw6rZgTBHw
vtR7pCwK31hUZVE+xHp6YDCRgoJjWGnt+nVxkHLh+b9XUKAN4TXKE7Mq7SG543eSjBq3wlZbPkY6
LMKCvZwvQkq6nj1jVZ8LAbFec0qJ6BbNL7riLUzsgy9bFg9E79RQYjFmXKMLbnr5mYEXHlfml+5a
30BKmQlpsVDC6C/591AIyoy4PRv3XotuKERs1D1CR98PJ2PUflA6vIOSSi3pzsRK1NnrbCqpMaU0
dI9sRGwZuWPGMYVwhGYRSdPcoI2x/lz7cf322LHcaEpLWerokvzZONmPCkuzboy/K1MA04ECDjSw
+lo/ObT85f4uQGu0tp2pcjSpcF4oXPZpC9mh3FgK6V7+Nh8NjJeEDo08VVjOr54E5YPcKq6U6kw0
2l8dj2Vy4u+LheTZx55NtxPzQqRSv54kzP9mHMTF0I2F8Nrz/uxGtrfy/N9kS0uZ4HggIYRmHKvf
yBn1vtYejL9YL+x+JKNZi+d9wQK6a/+cPSRBOt6gzckKOljIA2js7xCYAzpkIqsdVqka0jaGg3nY
2KvUZH36UyVQl8qv642h3SsLzUH84jjrnSlf9pFchBi99GVRHb/3YhCZyvmkcvgu/ncMh5bT0g5a
2GuKtiMb+cOtaf3HMrbpgqGirZVZm8YrQn6PwpF4JFiF86Co1Voy3fiFbrfq8g2E1jCqsHxDkC3T
KReLVQlhTIEgOACyBDEoOWno6lCdRbBaC9ZP2W/CPjlbT4BvbBClSG6PSpQhVR8Vlr00FFCw+g/V
hrtYK20EzXPuUguUeeJGsWZ2nTjum/1r8gUu+vU2TVmbpQeEZ8CtWm3tulo6h6+b2YWMJIUUnJWO
rg2oFEvXB6WftVxfBdzhPAWRAqGFcDshyD2sVQlNj2GdwpkSkdY3dvIw2UawP6BQycddRZ4uQMDM
wpCKmlshtRq+a79CqzTW31xgkQUeaDp/98tcJD8z66Q46dkDVphmVi+hzhXMawX8ez/ApKYR2S7T
WHmw3aVzDwwOREEDsAqs3HUysLDb49LJoSSii6cksB1EDGP93ijBNoINvsQj+jD3f+svNJHJdxTT
86bMCgorzX0FVPIzEm87tfK+MOcn5en3z/LXOxjgU7NW3RUnxeDU+tzWkV0IutTgWD1+PdVPgsck
l/tSZgNm6X2ypcwCKfhKEdh5ueas0af4xQhb1hje4swGasWVscm18JCEqCoFPibHN9UJ8A0grdLM
iLMhFp39/UwPMlYEC0DObGITGhXJcDZrQQF3oZ2K0ixXbjqr3ipZGtNkSeiwmJAZlSctWI4oL3Gr
D9qvbcJFBX+MVQ+nD+smkKH9b8KokD5dHfy+hHw4RVtc+JMdTqzeXyM3xK4CAyP5zeG4KImMJrJW
B0r4oYbfL+AaaIyWbNWqLhOC3R89xLqvBbEl5zL3HbYowP8rk/kPg4pubBpBHQo72VTiy8DbUqfR
uq3eDxtonIwH8UUTIo1p+Gz9NMITfBCjwfW8YPOLymJqo8dCyKAA/fAnT3cU+ARhc2TwFhz4tlsj
JFHZo16k18ZxyXqerirhJk62lTz8YIe+S0dgSjZHhrpyc9hWBAKzLVNGhFaEpCp6gSfoFBuHHbDZ
yq5uhC5PcELJ1661wUn/9Ho8CCEQw9pVIAEW9VahUm0oLGQWBfWsaIVFZEQfzTXbXrDOeEb8PjWJ
Fqa5M93mT3QAyo/+OUvqIvQDJuyGd1Y5a7WlyCiYyMN5lNIGwsO8xQj6d16zeaLdIn6RtWnPzJb+
iEn2LG6jYycm0GHNUHEzD5I6SlONIcgDhJDKw38JgGMeVUXC10ZBfW0L/h19j2uQNeWZyNJnNvNr
NJfkm5cJh7F4Fq/qmNJoo1Eh5AtMZ5eXomO7vPUXRj8ga8cZIKffywR/Jqixe+87qrl3SYQnv946
0fOP0QMGBAoOkLL5I4xw1ZtuEu3L53eTjL5b4AHb6DaXKHmt1sauTCpi42XPnENQDpc4xoxS1UWM
ebVcI/smRPAtwcEjOI631zpMusrUK8/rIrjVEsNahtvkX0gwHkrpRJhxdRKC09fgJ4hGm9qf3PbO
nCsQnB0QGbBhiIRpeunPW9dDPVgbdMuhoN+Gj3DrDpTf2ODnS2CM1LshJ1mLP1sy2ULNuieb21Km
m/SL84eJvTG0nzprrzDNmsUYdSkSSuEsrMHk8A+3exY31OijGcS220soZfQfcPiCblhVJOjWz6wI
4eDTpSX3/Z47xjqpEt+Mvpa67LDpR6ibfezhEWkAxfB2NUsuZJDsTaZwqjLKlyog1ckhRTrbu9GX
tOAMvJpUqybmHzZaXE7zRLhvEpQkISAWUtDQs9WU7xSgIXOXcTvnRDnOeGPcoYNjx0OXlZ69QwWe
BKZ8giCldImYrtizZzSvfexmkzfdvfG+murqCT8Q4kwH3tS/HFBFKVGcAdWkyRv/OkD+FliFgJmW
9ErRLN9dqng5C7SlyGF2s8v/OctNAT93zcUpJoDPt8vbNwnGwnOh/imGTdmkSPvI02a0w/bgncfG
mF6ApLSaaGTNlg0C+7fwjWhKRlN5Orm6ryAMybsn6Nfh4DPhbhQO/afqwPZjiaFQe2AgJKMJ5jbP
cCzj3n30mLW+2vPWvCYyPD61LWg3bDGk2Nic/06D0g4gusiFRl3M0YZreec9B3fQ90YEIz7jnRZ+
aKHylbtUCfAN9W0RHpqs6hzyc4tvLpuKEkKv9m1KVKgaU5lTbOrbyT1H547WdCgUCoJS37am841i
Uh72HUpDxh/xOF6XpJP6lb2RO9WwmMsx9ThO2RazrCVN8agl5k7tAk+ZwXiVRZKGVlR3XYjwCnVz
YEWheGicSPYZZyrt5isiXWFHwnKF/2v7S+IuyhL6QvRUz1eV0q3SHivVNCp9hUdQrkO+n4RRT8il
WS2Rqfat5ge6iUk+XFOaHHIOs59+m6LH6depobNoeGczAEPdkDXvsNY0uxkBuQGuLJ7Dra6mpUwc
Do/+OT2r1j7JQl8Ceg/gNiGgvpKzfLfLsW8lHu5fYylwCXTZCGXmdyF94SP/3CIVj50XXPxF13nS
i2o6N6sIMJcaCQZm+M4jZ2OutElrvIJVstJoQROyz8vfsazeLuhxBlKIs88FMHTD4vzFv4ZeHP14
K23C4eYeYNVnPReQN/9uDktTg9Fkg429lGjO3wXHoreEYjKuojJMBIdhfNZ5Yw+1+EKy6B5DgxgT
5G5wnfE4EE9GD3kSHxt/n8fH5RsfHQVEap8z4zLEKMHsmz6if9NbaxXiu1/vhjpJhFN+gmHYtaQx
Y7N/XMG4pxQjEWG+Eif1F/WxEdiXS0ImaDMdOScm3nt69U7t2y47pwnoXUm7pL/naSSiFxBm0OKY
gRfE1P3ZmosrLTL1KIZvf59atbPbCRdX1dRnThkzGTKBNzA1d7uQXEB2QarKCGqivHYbhkb7Itg5
ArPhYs33vLBzrKL5XTgJRq5sv/7U6MlYWeXOh5jjILqh/HCt2eHygMvjNRo9UfveSXwiXOeZ9kaR
tbxXvpjkK1tsF0pE7V48C6wJsEzlFTSZz256XwWNma1N28gR4hLTbStx+f68Tk0FuTy2tr5cPV7c
njGa4IE5dTuImRbFEAt1Y9QapkLmbtw782YZEqnhhkgQt+xQay5uqeAd/S1zwjx7ZpqZTpXH8MvX
fiJVJbXJzOEeLLYMQFGnFQw1WyBefgLCrYhlT4ue0vKglS2dzLyU2g85umi1PTWvEmqG0ud0nW7J
F9QXQh2pFgS+sSvsBL52oPeFnSYetp7XgdSobT6K/fVN/3Rc9dMCZZ/dBkgeSBp9GmG0phPFtuRm
s4YDKumiVmL6amFmj+eiwsG4RC9MsufNWkMQwllTgRvPcK3zNHzIUUqS5pfOfiAnVZQ3ji6cZKhW
5qyU9diKYiF2la0/ZefJHEAcP9g6ALUvMzuUzhIQFc64CNxO0zTx7OtHW6hA52qzAta7d3rrFm8i
UflNvuUrc3vYPsGReFj9aZhXvwvPXzigl+vJHflTM2GD4lL1L7u+tUHur4rBpfeMmxR3CKfheI+K
lxtIzdiS1Q8rVTNCCF9AS1hftjxYk7eiTYbVw3T8WaYk5l4NfeGmQ3x29h/x14TMmRteIZKVIEIh
Fjz6w4nxhwZQGe6HZaOcf8O4aaRp1QAX944S22zJpyJGYq8kdS16fAGNiVbm4E7xQ2RwzLqhRdk6
l5XLpQi1SBx7+8RmKiLA/SQOWAIzd8j2CXG+7s4X5kVYCi6EFUV2CMJDanunAecnyyJLDsYMFx0F
mRifAjVw/sLM1k0xeSrpbypU/rH3JMw+TKKxe4zuSv9HYY30I0taF2TQUaA0JV/gW8YQIDLzkQWA
Ls2IeBP676mpN12w3WZxiadCaLZyWGQv9PDoIpSYaJKiEquqZlZJCUXAJemLvY016zDaYOKZFfH+
zjoy7iKDwsP3jbKXYRkFUt+IPJHo4d1n2xPOeCXvloPtNBaPatsdRL2hr4hCN9RmfDTGUL0mZKWn
UGTbKAdeNzTmlMXbI1g8Nb5VUPx/2I6enDE9XrNUj7quyWN4sY2CHHg6sJvYzVkUX8G3ZemtHLTJ
KhUIYg5ah1KRt1txSHV/sG47gDjRa7nZL96YI788Z28kYsNlRQf2f3dLubgJzK9SongHCDMln6DH
ohPWTax1kxoi2QbmY8zRsxGWJDVwxcAbfz+NSBXwatF7IHzw50e1ecOQirnTIgVZXbtjLnYs9hg1
dZJ237y8wqTeSmL7LVoqh0RR2vY0CLY/au4ip6/cL2Bvqn5KrKBvm4ovAtGBHXb770jz544Icmq8
96zG5u7kwLTgKwmWGK9Tm9I93Vi0X/iRMrVhmAMQZFRzM8kDg0MePOpt8W8DmDWFJDzaq0T9+jkd
g3khGC+yy9lebNHOlfVwRotlTKD7Ssy2/0kl293mWnP0FXk4/ES8Z86nH5OuWAKzQum0P4DpJfy6
jfO4iI2UAw/VRUeNwF4W7bAx470+Ps0VBZl7ahJVs0fddy+KC5zZ1yTDu0ExWdLZ9aYIsFNBmyg/
PD2TZFLcmdr2WMNpNjK+Hfkl4D/PhK0HRrsXchFv7NBJynuYcu8mURqAGE0hu52wso8mjriwtRov
pEFCVPSiR1bL9Y1WcFmD74X07ZxS5K237LFwM4DOep9MYMX4JajW3XtqrKv+dJg69q3aV/+fdVu6
f+I6l6G0WlTtkaKMeqIZS+yYt3XqlwDCHPLQdZPvUsfV6/CjaY2FbISVDMmY/v/m4rBygxUrlqk3
yosP+JYQMgl2reslqHwQa3rLjo/Z66CMKd0/up1UnDmz1Nn2Ii7vT05TfgeO73s4Ph0Xq3XuXlav
IwhTJ5mIGxlE6kJRyKuYxPFrfNXhvRF5bmezjhVpw4Quvk7U2XY/pZeccUo0PU4ciJJAUHLb3Wva
m+Co+/A6bOM7jzOwjJcglMCQTKoeT74SZ4uEvuffV5YgcJH36Or8auk6fzqu+lRXF00lhCHr3JKj
LBtba4aX3YExYjTrHE62kFC+W69PgKGzAmU0c6+tCvKL8iuVFDE2KwZwhaUZBi4U0/VMhx6Y0bTX
nMYHbecKkKWUBVU262gMIZNXGmMqQhQuVU3Uw6nEVfnAo/oCozKE7WFBubqiJ/W9wvvDhL2ormKa
dj14HVxeCFeG1OyopB41DApNI1ZaTCKLonebdR/AZ75PWUIKBsCP3P4QRSkehWPvTiAWtFbpQ8De
kPcHkL6Eryrhqj+Q6SJolypBVTvn+AIHv86CsGbcBCWXs+iMqjezopiGQc0iUp/0Er2uAwLyaU5K
vEzwbgf6qMHVuGgAQoETU+YICSjmkprnHtaFKNkAoD7ZfvtgRIU4UuMASjVjq0i/qg8Dhjtt5ypy
zDtEObHgK3GSAEUL2eA2KmKRh+4Pvv6f+wbfKaHZgFbdow9MdGGQfxqe4a6+Dkh7tMHbHtVPGSGz
fZHgriGcIfxjk0xxEgM6h9nM319XXUTbBGoNOUzV8KG0XCzfylOebW23pfc50hS6ROk1A2tOxnZc
uIaDpjntIGi3ixenRAnjJDC5iTRZ7xPwuAzz24HmgNBd2XoZwT0G2UeJv8gu+r/9OAlD1vRAr7YY
jPJB20CAZZJx+IpATkNY8y+SrtClqpNFfHVk2jhSDEeiYDpatYbO2SgbrvHTYkelar+0ExMwFieI
EjM4n5nvEhYY5TWyTQm1FpL9A/gMFJXS79jAGoiZ1cePy3XmLqElcDdOJBmmyWeOg09LWoklBYbm
XJt0KtA649/mRJVLAlwhFw+XTNUkGgDBZ7CNzbHygWplpLhwF/OZZGQijaMiRxDsHOTrRAZB5jf9
XNcDeJI4fuIiygKr9WSBuaFflbQI1FFhOUkLzjZgVY1clg632EYX2wLyg1piWVeoPlKUxPvh07nJ
0bRe9wcqZWahVbBbDtQoF27zh15SKnsKGKua7WeD6XEDqaWAzsvQjqImH6/ydO7WrBU8lEvz+iRP
jTzlEkhz4xyEDcGHHLEHubgutrUTk9UCde+/z5/Y0hVGjELcyPXzmNuCTPmUeNn8DrwY5rc7RkLk
aQXWkL54dO2GxSXPV5mDHTqqEZz/O+5W4keKVF0JNID12hXBmQKK2o+tv62EBBMy7vmSmTtejgOk
Y+dV3o7VlKMMroU4xloJdWTOYDjjg2sDVlp7bTIdhkFFNmqQuqPc1ZhYhE2ZU0c7hDoCc+Yg04t/
eNYFGpNaELi4zK1SDurmkI+SbpRacGB49GN8fbnfjYJ9qpR0cEz1LDidgGG9yxwKOR4IPrROZOjM
LEdS439jauOPK7GpXcA9iHhCZcCJHu5qBZ/G8JJ3iDXSlqr8aJpci7QFCxBQfUOo+T7aJalpjr3z
8VMsBKg1K3jtpSEkgSXGkjxMrIYCFnwU6EhrGhvtOOWLKdcY2GAyo6BC+jlOGSlCJtyWHZ6uykJ9
xtOPq0myAJ5ymDRWuljuQZ/aj2MscToiNBnLh9Ltua4yc/MDGLoB8w2ejMcE+WcteT7g69izPu+X
6MeJwtQtb28usq9iX+0Ew3fpeWNZBQkjcv1KnqMzqz32XiBczPyF6VzA1qXEhf3VQ5DSdoL6HUub
yeCgdS5JRZ+y0j/s5xPH9FHR2L6x6rBWZSQ+v4lYbEvE/PqRLRpz5OcMIxVSL/2EOjAzYYbBcLTP
mCpT2BGCo7/LilZ8NfYbqczTUu07Wo7+8SSSe+Q5pzdqvSkIs8OfQ7DagzK3F68WHdyjVcSlH33K
+LRn2h9tgmQHZKgxlKJ3bGuGUvmfb1y6vXL24+NoF3+Gzwo2AuDSErMgT4BQ9GYRMS7CxaqFdojy
IYKGrHaTZOF5QJ2cfzxNsyAtZvRqGX5J3FSk2sKIC1JzdVj7ZnCqJ++TnYp5HOyab4P9Nwf2hj/A
njZCDQ4IYVhe4hr4uvI6nerJIoaf6q8OXnOzrfK1hU61sqPsPKOXWsR7V2kMdt8bB/W4bfxe6vrt
L1lSvTyo0MGcEpMXXMMhOGi1USk6lyJmrDe5GDnxuT1NKSpI9UG3j9dX1fX4r//LIEJNOsTz3urZ
3G7rqW0r+MrwL0DAtkgUSykVppv7KfeDlO61x08q3Izbxb0F0FQ8dRHEV1TqEw1DD57L3pD7TwYX
EVgoBM052j9WY1VS+HfVal9Wo/dU7ekufXDLnwwLN/RWPoRjrstT/s9zsp52zxDFyAphOYqvCdEU
qSwNQsN4+E3BL0jBEAnPV/FupfGriSWo/Wp6WiGVuIASkPd4BgntjpcquyFc/udRZ5FI5e1QPO8r
Vu8pzlxJBOeEc42cmw7XpM3lD3SU2CXNp4LJUgp9IhGzempllQFtmBNyh1Q7cMCFuNFc/xC/xHfL
WFWHLicN4mVQou2P0hauFVgGY8J9+cK/PDgZVShJJkOBNSH6sTqPOWIp9tWk9P0ruaaqpjMXRLh2
VAV/tW6vxC3KaccGEsx9C+Xz0cFX35BRLxI8fsufTJ03bncg8KPR+BLrb59QxjKLwIg29qNTNsJc
o0GD1MwFyFePoyKnR1wvStQ9y4j0E0ELW+E5bS9bW0RyenEtSV+6UBXJ/2roNDZ6ZzAd6GLGrtG6
qRxjDtfkcGxF8xpMxGwLzp/p20h32ERbrqYymfNjyQICt3gX0ZjHAunPeNpPDEMuTW5EGTEqt6uO
XXe3f0MQEMVfAZfET5iepNKtMcc7N6lfzE8LVS0zVFE20xv5d2h6fPqtFQ3fRRxysBbdpB0tJrNv
KiPch+gpBNRN3Dp+lTQMrmNjvx8j8+Ls1e9i3Di8C6nE/DEV3UDlTR+D5qSi4UV5IZKbAqODDQwV
KKDYe8VfK6cDsw75JJPJiiDdUEpnJzqoJlAd2blcv7eErA5e/RepP2b0/mkevuWNuJLztSSCrDAt
cuspQ0kRPRt0QBau92gmDewXwM2BblRsVTeHxGJ/2SPyzAD/vRhbRCXzlS4eIYuML9yBkfvk/qfN
ykhjaRVSCUXjD8k9p5uLis6ojFJ4Ji4RO5H8y0KMM5p9s2FSHCxquPpcQs4nBYY0GD62o+UVC5vT
ExMcYNnwn6WfrxRN5IGPz9/XD1k3mlNH6RHFT46HUogyAUUUWM19J/uld8aiwcIaTA8ezMAx1JRx
dFEZeIbbWzpxCLap+b5gBR/bGB6RpEHCvK087ESJfOgMcIFlVnDECK6DZJFkEpnb/7VVFmYY/Zl3
eGxvJU+GVhckDTEm++qg0gI3Y6NDWCUHf3cYSdjJhmqKQAM5yuBTd5CdqpgtOBCMgRXyIHDw4nX+
d9VNSbHkRwkeeg3RLTqa3PJ5omzZEk9gbWOLu5/nHYmCIf0378aGCCdJNYooDd8azsoV2ef4gXOD
Ffjxee0w0aTleAFy8pvfOK+DuDCtIyn09dYm44af/OnDBi9siYmjHvKQZ+x/9uCkhkWGybpxjJ7H
6Lx1fRTalCI5sXsYVZwKYO/0ij8TR3rRZxmQNo7FJSDfjW2A6tOuUwnLhhCDVt5Z7mMvgNlKXVDT
Maen77SoRKKGQ7BqmFxErLhCC0Un6YY0HhHbVa4I/2W20helHt6G7ziCd421wA/d2Wc11dAnsUF2
WCGRe20fmZPWfCnAcp6hbb7IDic040iSABJuVGzAebe/IJvQBKTePnCAqa2PXZUc1IfYVCWsJSeL
kLHR4yoUkieS1GybJamGxaq91lMFbm3XcuLhQ8ugjm2/gLFQ0YhuCFk9Xvc2cjaG+0hgXXyOWv8J
KsCmYr5mNCW7F/anbgTCoIWgStlZMps8id0B+JB8C9Wiq5v5lLwl5U9CdtqJUTnoB30mZBQT1iBE
UOSfQPJ5f/xOJTRLeLHYhbYEZctGvvXX0Iq9KYa2hPzsWYwnmwbw8DyWcYxCYFCj6m3AeAPs7WkK
8sTNtHfnyBqvQvJHWbAYmNzwkUYI1ooxyEZhtOotBLioqbl6atoT5Y01JUILmctSSGUmb2ONVf6C
nfI/gtnXXoZn07/SAYGWCiT1e2PyVRjR7RsawYdhw0mmQQTQ+bwSEDZYiN/LuZbEUstyy96MPioq
mmO6DGeQK0a+xM1aSEVvSU7RjkwsvwEzDL03dMvlWGg339A4RBao46CkAZJG5i5osMl6IkTL0HBP
LvoqZJOUmc4kDSq1nzMhcnzE7JN9I/oKrMB9PuISE6j0aEir0wSAwYXwGzptpaGKxkMYW8vDzf3h
0OG5mXr1NUElvHPLhYejhDfyuY2U6glKuATDuT5YwjFDXnlN1Nbn5jT/7G048bUc6yuqc5J5d66T
OaJJKp7JfpaoEHSo/jgDMLxWFL5bArkGC0mpwDDS6KYkPNjnIMcAyI8borI9OPCoCpytsFiHbHOi
A3mXCzQnrlqHoktJ5/xEWOR48SqdbwfJ5D1avWKOOjplEm4Hz88VZLd0f03vMXOw91DufJVf9aol
L/x4yORcBxgJWN2alV099teSzCnR2pPvHtorJBk51C2VlTys1y1/QmNT04ug1SNhy+4G9ev44WgD
RR/wgjqD/A8U+Au5CenRdJ9qFRwbD0cUpp4n4m28DcXtpy14AMYP6F/sBDlVzYhYyXcAol1vqxAJ
Y9k/DScOp/4AxLEk5e7/bYMCQyv7GLGmDBQiyVqBq06YeDfMv1JUfQ8T2KLc1PWrZlueSCoAQ9Nd
vrE5vGQr3X54aQQjWyrRrlpkmHrjPMdpwaRxZ6PuvwcP6yY8uATfngMDZgvLVxzTEiCYiiVF4PBV
ZyzFKilOn/9vTSa8d7k46YqNzSMnmznk8mWBcMlOO1Du6feGO8vmUvvwOdfYPVYjKsyXmIj0wVd5
kHh9FHxUkCTNAlVtg9FY2/RsDSthLuO4VOTAoqNMJmGJy2FJ0rCU8OsU070m0zUlZ2yK82FdTn8t
j8gQI9PJJL+8Hfcv4fF9zruCjBT9rJXYvLfIeiM/3qpPzMvTObzaBW7PeN0JF9Qh1pcEstwl6GBw
8qZ3QPC3vJfW69OlvV5nJLQWvmUXYAVUwkf1hgvrKMoNawnB02QcuUs0zo2soTsMN0uIhY15QD3G
qi5qAh02laYsBNYyuD7xEC/ZD/UbTd6eax7tSTpUU/PE9Tz5fuUimbvTiVOmpWNvZlkqlc59475u
ncBLQMnHtQRy7dWkGyxUqHzrE9Fcssych0FhATtFwh53+RyPxc3STop38vFfQfo8nuW1fl+N33A8
CuSOWoOxWRBMi46TPYuf1x0w01rMEM5VpK6RxZrpAAYqFkISafu2v7+tfHd3p5/ym1PZhw2JKNHi
NPOLtr22PcDlTJ5WwbfV1gAM8Z6Mc9Rn9uv+UxUfMRadINgdLDOlYVzlhH27CSpgjp8SvN57huRm
rNjKfy8JRgAlS02yLpxwyUDME4XTM0Z44+iQ+odMsNfz1mVdwwHsfDrKp9MWJOrmxqyQfMD2X6vQ
hilHWh9ZmOa39BwiT/0FNtqMMNKizeivWQfVlxS0l9c/2M5izt+LLB7+d0P6LILPyBgKern05etd
TcjRdRmv/uAx/IWpGQUYPDo4kn4ffTHjQvkp+6iricuFPLhlGy5b/l6wi8dbE62x2N5yeqJYkkKQ
RnUHeAICEkQ7vfxDVXiJLhq4F+ieRajNkVF72W/3fe264UFYC+FuyUKFPGtgbNNcaASYL6OdNVW0
aOJFtnCoBHjxEmt8OA0BBH3IMJNzG58072dzTeBSS8wZcXeSkaxOxZcNcIyvDpuYMvZACQrAiLZd
908sjQDpfpUzpINBAs4FDsY7YWmLCmNXXHSgehggMYhaWA4wLF/W4LEnwWlJTErtTQVynk5JUYhd
/yJjyzDLopgxSh22QzLmAzYfxYTPeWNCo4rQpivCT4Z3Kz5s0X2It+Vwynp090ItigevNlhYZ+FO
qKuH0u+5Ki4EeEvXcqXpDyR/P9LwGQyRRDeCS0Jf9JlxguV7Ulw5zz1ww94VFLlAlozWnd/4hJ5W
VcEYFF30Bytua90sPjUwnRmcViUdYnE1nKGAh+YEGTzhplOrIl+4w9gsJ6mV6mrh6Pm5YBpyN9SI
zaMHfOfMg5HH+oF2MH2O0G2TCJvvk97jqaqAUmkVimdNUysCnXpLc7lv2sGR0Zroo2mu0l+fJn0y
3hjo4dygKXmDSvGoEr/4jEJ9k6lp/AVgWq6fvw1o0NNIwdEX7Tiaop0+CcLDFq4Krps/u+kvJbNc
Dk5mUTf8LWpDKtmNEXs6EPnNZz8FZvxGQnYpssJKBgO1VYlVtX++kxyUWM9APJJzOUoKz4iRV7kK
NGJQjBW58NmZukHghUvbYGil9rGNZQV8ZRTncnjGYWh2fBdw7kstgAU/AZgLYmAejizU/E6+V7kp
5v5Izfb1ue0rD/otDUrf99CLm0KCrxG5JEJ+WFdqMaWD6a4Ix84a3JG9KaVl/agcNW8yGB2pvlJL
Adl1Q4vcbsXaEYSoJbj8x5xFGd3uEAylMzo1WI8gZcdNWRUt30bcpAsIveLQTzyfLKlAaoqM/6EJ
QKmG2RdNWaxRsiR5hsAacinAOc2fiGWh/cEKTlnqEws774KH3xisImw1wWXKDnNuKvNQMlJ4kkNq
mF3C+e86ONR7PV3Ywy44yHOmLC01JX5cpv7E72fiwOKs+eBRNyr44+SQWWY46On+npMfX0SH4rpQ
8Pn3O1nZlWz14TeNmSjJ+uU3DJrwKGRGCh/hUOnb2zWG99tPGCav81u5/9gpP/p4wxv0kHNJXEIV
+0cp+UTh5VPbc4JNx9rDVFIZK6F0POCMjCOQoA9n7ObUR4K+1aYrvT2fkkhVE9RCUXkVi8tqNODv
5axynR6w6D5lwi/udXHbWZp/RUBOABbNhYx2wxjoo+G2umNvLtAFrKro5RnEkSzylCIT/8HD2ITg
KLWCE4aT7WSHlmTzHA7hDo2SNmM4Rr5/E8LzGfCBBpGf9xiYfRoJ8rO+UFn1eOVOeWgOfPPsPnkd
TT85cuAAOOP5V8J/1HSQjUf30GEcXf17QOtPRAQdqYJHDoKjK7w4/a6Lag2Pu3GUyMk4R7tsWXtb
uLtQWzHvD0qnMPKdHwsBw+zdoKdsctdYPjYYSqf3SrSGt8hPkUkwEblGRf0ESq6Qx85ht6aQJx0W
iOgC9VBvHA4AE4+T99m6Ddu1cRU7dSZGCLUwKlKryC3UQd4i99IihFv6yU6IcHJg5rDXPrpnGQeb
U0esRnJ11pkVsTV6s4RF2W+mazcvM1q8YazjMVOAXu5D2EAYB1HMnO8WNRsav9bPGm1YhRxPPJcd
j0lj7gomYZaCSW9wtCwQVhehq/2tBngW3SpPhsot9WouSJ1NWqfrUpOGF+b0Y4wmStqQyjazEhBq
FjWEAD1Dxglnp57zhSsEcyVCp5nB+NraE7oLFy9x2PzLS2X2MxyYxETD9e979dnqze1UVOJzbrPK
lxbJNdjZdoyGk3E37dZGLwG4TR/IMQ1V2ytqAR02Q1GAaIhxskBsIkQF+DzVK+pStf2Cn5o6ZV0Y
Y+NvTyQfJMqd+DGPoAsHmKZi6cZi9vmCUkC2plWGH+jcJZMms6jeLhYYcRzZo/Iyr4EwFtWBM1wj
T57xc2EHI+6hfi1A17CSVAszk5Vatnvikh3coqJPIf1KrZNMLa/GLK9cgaIoEb2+3c5GL26cK6F8
+9vGldXZAk0+Xt9gc4LnzmP+m5sEYshZoQKixzi65eht2saEuQ00+1F3SiZVvvJcR3r3M1a6ud5G
BYT8LeVAcoPpMQbZaNXO76foXcWBJVuEcg0Md06epQ3mGQto7+QdO5UHHiACChurhx8j8QyBY6T0
bNVByMAM178NoVT45+qJcwDIa4ZC4nJFkJpPasijnHdf6dv2YQZi5TkyajJ0wKQMj5rhMVubZcnZ
QEEfS9viAhDQSG2lZCkawF1vMRzCC+MhmyS0FcyLc8UyUmvkzmAp4gwSnWLz1CGLcPONCgierBEw
ShEi6C33QaT1686Yc+IcYbsPPVC6FmOeBoh27NscPJVVTFiPdMdpHLD1vwhJcMkNGO1LAbDlCRxk
DyIMQl9g6Bt1WpQSXBcgKtH8TO0r8jGxq7uk9J52CX2KGfW2rxBg35cDMY+AvCTKiIMNb4NtphZ2
XSkeMGTROa+Ajxb046UvN/Rr8MGrJK04y7qSuiq1uyT92ptSzYlsT+pHdpmFD6Ro10wEzT70Iy8d
3+rAz7ImeUnw6Cz5sVTdyxuZ7Iw4HukQhC3GwaheUswSJb0JZYwJe1xGvtU2ByvEph0KN/Q1JSyl
oony3N067wY9cfpl0vOrS3D+BSGsuxufYu62cG6Y2ZPIn+kZdmyc4mlT0iPAzlQMCCGzaYfBr8ZT
dTrmGUPLWmqjSEdWfiseRZ0jqvU+bjO2PbxanP4eRWtGqe9mbKqnKkPKJRyCiYp1uSIuuu43U+kV
I3O/uPKeflrEDVQjtIWRdQm0EYxBW3+M8FEUpbO6nEOqdKTcERkXRnJ4pmEFHun5xvkc9eQgMxAv
Cod6PGzTj5EWpg5ZNqQAZzW+FAgeh8eiUu7SPwqCOLzYS9nSoj/yXZlGqUUyEG4n2b6MxQv1Z+EX
Evg3mVzYhI43pWA+PefKxfxYJedeIQGtpDB/dpugylF41IDfH8WW9vFaatr/ufaVTpkyVz0ltHsB
2EnANQkiGZEmVCXCEufhNw37oSEPEYsGgj915gTSCl6cEqEEZ59qCyU6+MflFeBqkru03l3oK/Bc
ePWH3kl8XukM89sTt3eaHiwVTV2Vh669X8OIFrx5NhMAKcconK01f6YQnb3RKfcs69mUyAQntlCq
r9NBX3l22yo7LhyeTGqy5Sc1SMseIQyEqL8qq8tWFekb5GMhckMsdypDtfP7hHyxnkpDX8Mn/S6C
xJVEIXBGounLHlml32qkQvtHGw1ISy09oSTLBE0Ti772UbA4xJvTwyBqt2kLhOTiCjX1bfU2bPPt
e3v1QuT1GJgDIecgerk3hn+f1xN2nEy+DBzuNYgeBHxYvzKINRg5Yc64GqkIYXHdmAfi4bUugF5a
/ATvMM+RzhfQSNOj/lEOQY++vkHiQceanvb6jyGOeBjvP+lobOHBoXCcMLJFaQcbarZNLR/Ihu+j
MctwEXKqJzc4a0ivjGDMPgkO9iP1VRcq4Paf8G+GZ5FYZIS7iaE/IOLLXjA0HUGd3JtBOk6YBpDX
Q6vNElZoMeHv1Ogff1l4DFu+lqpXXhTYyUXiVI8p2i/TFXIBtR2fOtWAWRagUvIclXQzj4Ql2FNx
g3c4lQmpiSSqzXY26HF8JoXajrhhxfzp6cHKCKq1s/al8V8aDoVQYzUjNV6swc8SeERI4iWrT4Rn
MOd8tyqwBxVD0O22gCtmRJ8lL/BNgPXFlZFGg3u/8dk3pRyctSB+5OaJQ/QAOM7TtiUbHckrLgvz
TYWdwKK3UpWHYbLObSdjy34hllzRWQKTouFeJUtkTT6lKK5OBngO2XuSRvExrOcWPzg1K8UBdCIr
ra5Onhe759NrcCPi6NWf8b8JDKUnZhsEzdzjbp25Sz7dEhPHfE7sK5MBVik+gtc2aFVC4KHBJrfk
RmtJKPCijU/RV/t7o0J95jC+bh8mffENktbVACJz+dNqjtbltdNeJhgYOr7gTxPyLRN9q+Pcc03K
5yqq3RYws+T6R5z94z1XIVq9a6EwH/yeMS5IfFVHYVd5Pts2dQM1g/UU6phXXjuekCWTN9zAhYRw
ZpcRB7HVVsic1udBfpvMsZB0xYInLp3MsXXCW+iB/Pzg4+YM3n9IJQU/mKITSHoYpngP5oppXDru
RMktECfT2jtt4dEQ+hkHsgrW7ooFLiB/ARMdDL/0lD6+bfL0aOOqf++bbztwoHkiyD9bZVverEgP
tPzwAWtymsy7rqJylJD7YREecWLpHb4gP1B9Y+JIOmvq8TUfdOVQr2XdBSX6r8xDTuLsv2LUrCo1
X158p2IamuL2qslcnST9N1XuSRFz8V153zDaI7koQrQ++CPTd5m1WXcMoNKRhywNNCMqRq7Syp9E
xlo5BKnk7TSHEmc5NSX2127O1mO7hfeIvwC5gmE45F87NHHYsYCd3Ay1d1oYjl3sgikxeduMGovm
b22W8tzNv1FbvQYsDcIg6TMP3p4U4i4iazwq4Gvqcmk6JmC8zdG9HLHjdVIuLR73p1dLzonTqjyq
6HkdiLOy6I5yB3fSBpzDJ5QfUwQ8gZTbk7G3t5b8lCW1ucAQy4u1QCcRtDYs9vXppnEcTl4O7z+x
8gSAmtccW5BYpJAPWXmeiyMbQwrc00HqZ97zbPdl24I0PEMzZAw5Cv/Dsgn9I5csd2OwL10zzXwq
sNbvmtL6EX8LIXeo1OsRac5l551Ez9m1D+tDRBbXlFns4CtpL79+KCuYdJY2VKwrEZSJNN/xqfiH
ZVQbB0JOm7dW+WWONphhO87hHpwWLmdw6MErD3/XAHjrJdMTeIJ0y7WTx+whSgCit7LQLSzcSCXh
TdwkXg+tVe+2pwPSOEREzq5y821qjaw9uHej0CuM/80LN4Bpnvd0oH21yXuXld3tgco2Hgt3BBXE
du4+eG/o4M/lUk2jj1z5bWuJcTNG3rt+gTB4Y/6Cbe/a8ajtIeFIiwO9jrRc4APLGgAdbDkgUMce
5uG2CXvS6BY64GvF+ACUoB/49nldc/TnxoXz1KjY98rmK5yqdbp3rNmTpRl0EtdCBn5a0+mr/9Xd
zWQZVGoZw5paaIW118HrJPjLXVuCoRPBRvB6eWx0xvwMOJSfDZQEj1ph8ntr5+wjGb5O+PUgVNJ8
PwMSUf60o+yn54ZCHTToR4IMqWzefxSdnC3XvrOXKqTd8C22L7MX6auVgaHtsDM8XR1kjsDvXIlf
pKwe30coCpWP2MSu2MT9COcfS9LIGXKbRL7j2DOe89EntYq5ANQgxcJiQrTqlJpQ8uQ4v/RGYU2U
Bbpeuotm9f8AGYi0jg0HGd/+SKd2IKEcBSXYqaxok/7tNS/vtSIeNSn++BFEIm3MQhmIi+6bPUIO
I6sZ2NdX3ux5w6a2vZ18Th9Z8YbcaaSBXmPVUXNdQ/9BuclW2jjUvenb0K699l3tI3x8dYmDLrMF
odrdYKiuHcynAtHwUOgO9BbDhwfvFpmiCaMRHuwkPR5OTLGiNE8rBcCHd+wGJ0MVLpkbFlx8Utmb
idSajIaoZQNkFBn5/VXEjDBMHyEOE9koYTDlo4yJKNZ3CYNFh7SQMzp/ZScHdS5HpQCqwLA9oYEl
O+YV7eHGmb6OdhgSRpkRN6bOETTtLssQZngMepsR+CMMHUIF5wUeVsPG4jJevu+Kuh9CHXWCGyUx
IHgkNTkztOkvIhkYaGpAfE4EaGofPGjL+1qJscpfJShndJ+5Afqf9XCVhv86HLvh6ZUskEOBYCky
W6ncJllTkUQqPhM9CnJC0jdJr3GcSNJyHjeRf/mI5glgLPY54SBHT5xcJHIaOpvuKkLmxuZ++FNg
wch+O7QG68NF9SmZCic6DpBC+2epU84VpERbufnHc4ZrLwYrJJbIwNzhD2pxrL9OeDXZE6gKlGpt
WpkuPieMQ+jbKIkdnTIXtsBZTyKyCwl2/UqpK4j74U925B7u6wDq5rnIe3WL7ipBkO20Ay8C34pj
OU4vdXSqSUXYb+7hakj8+lJbJCybAlkLEECllo+uaxoLidXE6Z661FAugWS7pleB7EB8h+iCGw1G
I275XVJPXEb1/acZ733VmdDmjbVPuvusEJKf9ijJH+98BF1hx3780VXasf6/nR/4MSmFNOisTB+k
V0em4vW6EUadTE7iQ9keyRW8zyS1SYkhj5CoU5YSR0Z643qi0z/omWslhJ6gJ+CyEwIDDQ/2ot7+
7TJVjU2UU9RpwXJzOnm3H8mA4TPU+r3DuM9SFuqG2ao8/Z3uGEQzbA/5llZvxqr7mCrNyEV7Fza0
zCXjqSFdtePLpVbWF06ylbU1wFIyknWfy2WprJUlN/sOpSPmbkE7BU538gqyp6SZbns77jqziXB2
V6SQgmTOVNk5x4/rSVj/CUYTN2kbQV7tODO1RKqTWday3UASBYRvu2IFv4FarsLxpbbVZUu83eIB
TKqcYQHyKdi2lBMdTLpcdyYLv4L8qaGdiSOsFR2za2wGTVAkKfeJEXQFlWY3ieG8eyvoEf9wKS50
pKmkA69O9CH/ox2plbbgfjOEqkouBkUIf0y5KOrOivgnx+dylPowiwBX0t9D4VE1RlB1hZ6rhwAb
P/RKNjqkqWO8Y+KRlQXXdN+1J92Ngnv9oj4m2KTOKp4gewlu8L8E2GvuRm2XHqoEUxBoiUimxHSz
t+PChcNY96o9OvXejy+YCWo5Q2hLYnNGxi4087vgvzjmgOeU4zs8ycMBQCCfHWlyCf4uiikjn3Ck
YZ/P3LYIBf6EjGubx+Mhn/LYn00SBJleRsgYP5BxhST9EEaJjCs83hMn54yRmUDSYdt1vp11nzlb
4saVk+d0493PbBeUvh6SAq3dFWip8Gqadjw81JXHhLLnATkpPjVNNhOTdHaLLHC6r1YXxI++WvUH
Y6jVtNFujBEiYn5y8YNMHet13abWdlWCNBwlFqWgNPGx97GZP2JN3itOK8yQOqqVI+zP/r6WhTEi
tn4UPjlVXYkRZq2UZzIZjjdcbVvVKoMvS96A5+V2NsNXfWHT7Y8WfUf6llzLpCxYmYR1UZYB2IvY
DBIkdgHlmjsJy+P8gK5O+pVBTcPT4sr5AZ9LMUVfgfhKHQ4I86CCwppsmRohBT/22m+4Uh4w3QXW
qHEh1HFvQWKGvYO1z942R6ecljlhciF7vDRu3FXsr62Jo8JDSokvrWNrnRbMpsmidsKASGM25NRy
WPu4IA0HJfabXOSWLXz+dzRa9179dcI9JufrTO0eNZ+92M+jVLNqSPHWlziDrHkX7pC8gCZz0pnZ
qhaTXRIWn0hnXYEvqXUPiCzKsUfoCHU0g8t3XL9d5A3Ltcnij60fsAZ9deQ5ixs3j1qu9vY1faxA
mLg7QZgdrE7v73739kwvM82K717Efnkag9uA3MGlXBhX+UPd/6QdadNqzJ64qX4jA1IdReh3FP/6
rsNuLcZxqzcdzrRqQ6GvGl4WUSj05t4nmIaNraP5PfBYlXrbp3fFEWSp4udJX0vVeFogNq+KeiHW
2zDvrIXr4wc3htHVr2FgXBllPjokV7f15rTP59zJnvA+6mjvqZELSkHehdpGaCeIQ2EVqqF2JyZZ
/42k923E+OZXHDPRVPndqNHrwO1LYEBI+2bSTw3Ntg1rLfs4B7KotyGLdo1uvJxA1YkYYXEnBuJm
AOPwc+JqJ+myMna967+bwMkey7NrRJ6xKbRkdvPfQNhQYliknjcmRC6KVJFE12aULNX5zqsNZJ1m
ygWdlDdRiOkCAFTmomKdufvTABhCSAmEioBl2+d/wyq3L+MoaQbKoEyKYHvJaD9MYi43S/bPqP4E
sUTA+czgb7POK4OUBGwzFGg9KpshSTQiqABIydeHgB96kg57hudH823H6+2ZJ+4La8M+8kFDll6J
ebr3qNzvaBgDSoocd7D8cxJIZdVBomWqOdgiOEPpw1e8yk/PNKylR9ZTaxHOb98yzpN/uk3BNdNg
XiwdcPPD1CHH8+SDStT8hxYDjJBMLwhlFhFEo91+SjUlE5KF6agVXNkQP9ldDdycWvnUwznWwTZ/
orwRRzj6F+QjrWofayPWZ+Bt2D1kffU+YvIh44Y3Gxdrcs70btg3qe26PO32rRwOW3XOHbIu9JP+
OtstTdiAE18MfEgFr3gp4iI2ZABvkwmJQ143/ErBXXAFWoXlcFBMw5lo/cFwYAj41zvmCQplrcO8
LKv473/UCkOw4DnMzVvc6bWl75dhPtJkS8RXtL0SaSpVfU2nACMzThvNN99ZR+QuW94MExNHWwRL
BFO5+kXjG8zbHPNzPNBnXDodGAuz8ifcpIJrIKdEMuiqbDI5lMqTRUivcRn1NgT7rbeQNHDx8CF9
p9z9wFBXb4GZb6omYJ/+4nJrbr4GcaTqGIulQ0viJD6tiu6SLCCwbXq4NBtdzf+pi/0oVoq1gzIi
G3GXmruAyy2XcjOU0JuXf7vRN/MCOWvNGfioqs+MFckiXSIakf1SCcToR2pcUnRa5n2vW0KnSECZ
uQj7TX6eWTWrXysOFObayNv2Q+WOPHvaVUb6yT+THX5Bd//hxL7wUEYo6Dt3G/QjD8idVo5eIVxh
pG0FhUZPock06FF2roWrRsetHCOBnE6uhCj1DInRPJquNfiZ0JhP4B/W4D+uvd00Fs//oBl4Wcjw
OphKqxZJST5LNIv+lCyBQvd6g+FYzDWTZhCozk5ppECEPtjWbHoeDVwudgkvRTUtKyR36PUw5TzJ
GNvILNEC6knbyLsoxSI15SferT5OKjxYQ6OPm0N1qyX5y0ETNeGu3qjnfvlK6tEhVTHLHEGqWkev
ZcFsU0n4y9zdZKj0j66WKMNH1knPsUKjLAyxZjEe1NUEnn5vnwv7zNf0F8vHmIVAqF9zHmzTC3Y+
QtuBQi9zXqXoecYnnig2NxpMuMxCNMlEwfqUIqlN+KVqbNX4xKD4KDsdSBwLtGP4nkIJmEDa7lTI
kbukd+I3RzGR/3NOUwOygGhVdm7IT4E47iKQnGhHJP2kmCNDzPmIcrEWgpGHlfDiUMArgS7VOk/m
Bn3rL2Tnebye7q2/FcsJDUci+BQKVavH7TvlkB0F4wyeosvmW/3KgoykPa773hwZVMVP6Ov05h6g
tPYAiwbdUsWPUVxcbT0jWJAZOi7tXwVLxGEQDnBHOBLBqsF6/xJg1Q1MRoDcc/3JVrxtHo2S9Vxu
AkRBeErjeSnSnlPGfc6X/eVi0sGo9AIaButwDMFDEImg+T1xYIAubYJrug5yp0LHNlnHqbcFtgUy
0qbB/i8igavO63uHPu8zwaHHbAmgvZTmkeT2icZX/XBlZoy58+6doHWcrJ8RSWY+Y5NlTwZ2Dwx1
taLaC2jiqChm96KQWSJ+YbRc3TlI+gCGM9aKhc8YUXAUjoXXVqaKvczR3EjZNUeijMVPEU2VnVl0
5jDM2eNGAr95/ZbyAuGjv3ZW7TqPUIYHaPOloblViZ1exAterrW/rRjJxLmpFUWPODP9+Jr/a2hT
JRWqERzppWI894qTLuhjGac8Myc1+sEauy8fNXlqAtHWIEJ1r5Iu5GI2n1rABMe92x9xnvuH5dkL
c4xM2puaP75KBKwxhz/NvfkZgsm/MXwTYQqLEscDaML4jEhMomvGmPimlpLN83u/bb5h9HEbDg3R
CYAL3cuT2OT9h6rnBCOxLorGIF8qfNhTnXL9iv+EhHRrYCPMdjmjY9z9DIYrsJcgJFuCLAxDxxCO
DFsEHdi8YB+g2dtibegCPxEWW5HHL7HPKCFwCjXeFi8UYpZ0FsjeFydkXGfgDG+NYgZiThmohcFG
Zj5bai6dxYXwPleXiWuXgslPrN9T9wis4GO5OJjBO0FZaKm10zbnUMIbWb2dZyApmEBy/61TKKxH
ZqmvS7zwiMeqaPXToozbVAh5DOKo2CTr+gwv35Lc9SED383FJoKrHtAwfOFZJIRGbFeUyr6c7oH6
0fsYNfydiTTdQ3dvoDyHY8k4Jt1OHQzxijLz1brOYNW/pAQZO2pD8XDYd6aZfYNauTAd40uPJeXf
jb0dv9JCLjKmWIbiLSJdZLTxC1di4X6TOYKdHWxBbEm4nQQYG149A8nZMRguNT+08I0Drb04EmWG
BUbem2I7d3f7bh/tIAnItXQNi7T85RAyzkUdkRs3lQ+HstHO8E+oTxW7CJlEqAsELo1uSvwwouWL
AKHbDKes4mSchvWEtBuCFRgPyUa1IcOu9eEYgz4KbEE8sUC/4aWzlKgbg25kItuLTurfg/6YeNdZ
HnYhk9tWQ2iLmpdTKThBo3fB2eEKwvikUSEIxMPaWL3wDP0eFMz8RnIw/G82GMwLcI7t9OrozCOp
z3x4zYIzl3msF4AEdXMFJof+pk3fSAZa2pVVUz9AS3gU4KjZtdLYurxBWusftmJCPTsPIZih/nJE
J2ZXthA1TrTUI/rkzZsEV9MpORHaIRgwvExI7C5rvQ8U4cqpkY/rrQ/HoAhFVb3pGyRBz7fRKQRT
51RZ+phs05KVAq0QkJYzbwVGGYXG5OoKXs/spxe+ZjLp//W0yc7+xREDad5OTcjTp5oLZs0rzbxC
f3l3rSWdm1KEypbB0KCpMZLyKSHVmiFhKLQddhlVK2MWI8pqClYLeRgA7XshdrREBiwtEp+WZoRw
bFPtEz0SF6Veg3rrlRor1vgIBLKARJa5JpgQYMlLwe1APivBOrMK9lNocB4c0Wd78G9aMV4biFoG
3KpMfjk4P0XGadrxHoYmYRtC8TZzCLjt3aMh60aa5ui5ELbwMWAv1LgguXzLRM6sn033B5tj2iBc
4ZGCXLMSo/S2bUmR3lEF9e65kNV5TMCr+FH2YtkqePai7x7IMKKoV8Dp17hMCgFVngfhJG/LwCY6
elF232V5LFZCSMX8Dttm3Ze5hcPSxfJJRTBqjl0XmK++WQNCu/WQgobD9RyhzZbG1TfuCP2U3oBH
ajwMws++Xm6FESkmOJsVHI+Swby+26Lqog8nOe3iaT8vp3FfoZS+xWCzt5Il8ZlGL4bw4S4lxZNk
syUo62Jha4CjBiYDkpYsU2Gi5qFNtDZ39ssYMpdaz97FA06AaHy7SW5OPv73sIz4s4vAm3PvN+5z
OR9M1hPkyCLdta99vmHyAXa9XRXeu48Wymwa08v17igbiO7pTmmWioBMXyUad7RS5For9sfGbjEs
cbOR+1aolmR+Gf38d5rmYJxQ/DcEUDuEmvHUVe08FO52tzC3BP71PMDQS4WZRTxgig26N9uwT78V
X7LIOMdPNuybtJ3QyNosusVyLi74KQJQJ6QswipnfbDFK+t+tdgnr9cUqaWMa1qLoClTyGaCmoPP
fBEns+Kc2lXnshnEYeKArPw7o5jiqiKWZyyWTcDOdk8R2qA/4rhR+lCXMU+9p8/oa9GuY+Biifxi
HS7BmRT/11+hpm5WgBA90N/Em7XvruDfV7Ub30CbmpsEay5y3SHa/jW9Leel8SBWfkTFxcW1QtYy
g1lXx6K6cmEP+EOzu3FycgR/9gMrqVtUksOxZiEfEFCKvLR+5LBUtgvexwt62pbSCUS+6cs7z/WO
VDs/MRA3iBwk64+u6UgdTvBl4mwkPvN4ZvkbUsBIZTKtcRvrep8M1vbaezeH3TzqZE0I/AqdCaOP
I1VZLYmq5e6MCXgo2jnRBy8EONvVL/LLP8hYxXZk+yVVZAhGvU1SSRM0cps2qKQ1FISOC74UeAja
rAnuynRcKGOtzHbsUsRqBzlaSau/ub8GmWdfz7Ppbz29yhWauGZdQuQmO72upHvH0mSxiHkjiitt
6e2NpOXi8ANqnMR5p8Xu7HHe4fMlU9JySkQCb3SYXMrniqm1E+gaUNtDa6Kd+SnYg9yKuJws/bdA
dvpVfUZEl9ylbmcfyLAK2pRnzKOgRywAxdluRKd+GfOpKMWbACDdEW7VAVJ2xjSVIjO/LHctBXs0
1zPk414KVQrfRmkTKejQyoe5WCNQupic8p9F/LpdSeYHP+DmdOdwVrp+xOOivied5atweYJ/t+QK
NUwdoGkA4nU5A5RSr9K+Mj0nY8+PSmvzTjIuLm/iFQvYi9NYIf4ZRMQGQDpaFkAqWRepp5+KqUt3
GKwpTqpkqgT1OcI2zzazmA37O1E/wX4zMxzJacy03Oxnt6eNCDxac6IEJOP6UzHRmXZUAk9O4M8Z
aRPsH1/E30Wwqvi5DWyDjIqBqc8Ug4Z0Dm9+QRSTC/ForKzHxCciPtK+1Ucw36exggwZ0oXZquXA
UZ5mjqB9Nd7t1YD+F8QpUjARXpOh2iBH0D0d5ZUck7olEEGu2uop0uYhjQxexLPY4GAe5XEbiYW8
cCTNkfEtB2hVl6g/hYbQTNH5nyqy4zY6kj2lHLGOXtZffwyS1OOoq5EQV7+j3iZF/MNkkFWXLbQP
ejx+gsVnWMeoApUmaJdEMfccBt8PEWhwjHXZg+afwanbo5MDGT3kO1RlZxC8seX1burqUeGD+v7F
5rJSmadwpylMrGnIS8BkiiB5R/5xd7PaoZPG7Q4rGS5x0JqM4LN7w0DQAtJVvEiq9iyLW0Mt4nI6
CkIMi/pfc3qzCmHHJaz1y50DWBN4Ouad1LX7ycim/g+QXhGCLJiMHJNYc3JhnICQj1H4T2puImUd
UYsSkGbtoFCS1+A/Di2T/QKNBpi+JhjAWa9psHtLPwxNhLAJt740stMhDwWceNTLlGbFt/vb5CG+
zVUKvQ7QPuTqUox6VzoLuOGpz8+ooPUISW5BLM4BxqBSMzJ81gWj+AHJLZqv5NTADLW+jd6RGaQ3
v2j1vgLDWN+GpIyQpe8fbp/RTYW4UFvwSfwTHOM2zT4knyt21g1WUz4c+KYrlHlZnhdeZzlEJJ8/
F9i7EoAbbvZZSRsBkLp2mjFUsSpYTfZNLnSV3bnFNG9q0sFtl7zvCOalo80mvC5mwLiPbu90VlIA
TmJrGnea8vuWTksutz7/JzFm71aExE4gjUw19EGSSL6WqFkUK7NQeYaof9+a1wOyRtZQu1tzIg94
Zimz8dvrVvbe1x7NHaXgG3G3yOS4YoJB43tpZyVvOL1nSNGPP9C1Tjo0pN1FdkdLP6PYVJOdHods
i5jC/MLXEdhfS9ejnvr83czpgnU3EsJBE0lnkCt9gPDS3h1iK3/PnkDsFnNBsjs3nUDDABgVuPFE
TjZuFBh1lcR2T1yMcKKvqBaD84X6lXj5U5ISrKMSXza0caNgXwclwq1qrYBgOcT1LhgQVeNmSLEh
4GLhQpKlBpSkVc3RN86/ZijqBkNM3srlG4COWLcJYB9c1I2TbQPIVymJ5hhJ9EVwnFpm4jPGxlXo
P8zn7bGuJJrfzusZh5hkkoHi8g5i7KXgYhIi1DJiokFTrRztvwyTMnQd6eQ7SK4PgBE8r1vNvnkR
GwatuH1LtaTgQ8oyAp9A2KW4pO5uJ7nsbNzhELi9cZvbhKR46FI/35pF3R3A1Gvv7y31RsvysGlw
j46l6UcsQDxTeaF1/PhO4DO3Kbj6UfZ2LSjnewfRBYxKvPkAU+yRx6M4PnkLxhBJFvggDm/FmMje
ZMPCsDO2GUO1wDsMAhlAWduYiT8J+I/BCyeM8h+QEG06ZTwzKY1v5509rKzw3GNUg25++AOrKYr7
Mq1HyTTWiC+GM2LvG3HQ3SLfDvqvyvg8Bc2V9Z/M0pkGwaY7S6tVWV6CCIdP5uII0NcvheK3ud/B
XiC7rbcZuFqhF7j5R8CTzPusu2O63WSIh3VS2VPrEOXjGtUiIJTfL82rCHEYlRatDCHIDmT8KnXD
OTHFuaqtxqtCjdQEw/DVMdZp0wj91tomqOmG4Bu5KX82d+u4l5EDUoMFH0nY68rnoTkwShEZ5136
4AqW9DDuV47Q7R+rP7uwwUcgGvjUX/rzxGmf8eumdbE46cs44CrfXkJ49lqZtKao7kaoaY7x/nEA
jGn9DJbhQJIRiaXXOIYzugoz/8q9lBVTeU2Kp+pWUUuFEtfEV0Upm2eGxM+RddzVNfPtB11ezPdY
QZYYgGi88eGXIu9Sn/hV+rkVWf+GIXuVptF+BSrKdRUGP8L4NfWfMk8JSuVSr1hs24FRAJNY0MCw
mM8iWVjz07Cj8xGWTXVnIXhCpuQEqQFiQvkzAVK0oBDLE+RiSzcl84TtorE159eIE6O0YGcs2nXy
tFA4HF0kg+iJbEej5Jv9gPtYulu3jYIP53IgKyZkN3vJtf6DEdsbnNjT8O+UeD62jYUcy+AXn9kx
5tFCQ0bYmSMDfVuQ3mqLJLCSw8CkT17ZjdnOmicCOUZNxSLg1NYTrC7th0Oa5NTYheSbOlBSzvwO
K5xzrOpBAZLpjO7I82Zfcmfmq84Pt5eq5E6GE2RyFupSba/nZ8Pu9Fu9yhmiF/RB8zbI6mtGJ5RK
HjpNwAOamcWRr4LjtMv9m+7tc0LenTYmUR+oNKrKU5Bh5Qinbd7cx8Z3nhmrkZNqK7/PFv173l3a
185M8LyAa4DuU+SpybKZQPbl9pXEinQRiF2P85J3HXmA9H1A60juSouLJNZIK0CKvH/B9r+yy84j
cMUYGvYcLQbLbfDU2EAVg4XixyFEDns3B/Ngd5C+GPqgvvxocI5hlPPsHLFb2pTVtuFlcKtD0jR/
KaG31D1edrPdMKdMcYiYl6OKSO+afB6Z+5WxxHtxlmaDlX8d+Auv3OZpFe1TnR9nO+gv1wYfyAkJ
RDDWldoBph7vzEn+Uqpdh+5TfHTcHIw6IUYpJs5N+DFoKSLCGS9M9LQT0MRbzkRnwtoiD2sUu5Zi
UlltqBsTFrQy863G3O+qWzmz04NUwtgM4GW86sPXBHw5YSCaKDwiGdNde98igmb/0dNkYAq1Rjfi
2/PcF4N3LsaW8/7p+6mbqEbywJFum3TQEA2oBkGmujwFUzEh4b314CgnyWUnOzOiaYVyo3en08tH
nBw7if6hufTb0cNSu2Zlx47jPLtZzMzDSQOhBT6Km3WaaO0dpwoPgJBxyKCVoccr92cz3By1tPQy
4FXXxpQtvZcRfxEeS4cO7pFNlXS0aF9KVia8Ei/A5XaKGd/05Iab3kLi+dX86bI0BAkoqiA3XzkG
/oqnshQCEcUso8hXD4KokXuYytJn9qTnwc/a469QSjdnKiLNqY7OqyMWGt+ujHdJPFBdRHaHargC
mmkkUlSC3OwDEA+37qJsibwS+8U9goqfc1bYniSPaK9H11jtVNQAGzot0g9UJ8dPwFN2SFumgJSl
Xg5LrZ/MYNqnGOVpNwxiVYoXZk8y15ibeujvu1BLh97R1fzpu6sJCxlQSGRapxcPnVhMdsFJfRkf
YMCS8bkAP/wIjFEevObxnYWk91Dq7x/KhYoEdE42FKb6IZjoDNTI59kdoqTl7AM0RdZ5CJaPhE3F
bvum3/LOT9T+MxBhJk6PaGYqEeyGKV5l/bppr2OwTcLEdPCwnbpI9JK3r2jbUSdkxQceBv0MKSQH
d/tC2Fls1/NFW3f5MIJYz1+1MQw6fECZ9z52p/5KCvUc3C+H/lvdj1aLXaAXyVnuYMw4eqkeuP3G
5s+Bmf909XXLnXlS67bTwwwtGuRzjY4Qkclme7Njr98YKLks7U847jMBENzTqiiU4uqCA57UbAm+
/MB7vDF9R0ImndA+uVBcykvVE6qhH9C7s4gy2RjaeC20uaiFjEtnAtEdYE1K8uahoWUaxPIbtLBH
DDTrKgkmy9N94ranSlL9EPKMM3qSEF59Hvvtt8OOnrBtxC+RsMxG9GddUNLiCAp900yYQzT4LfN/
3tuqZ8spuFp686piioi2WHbVxhWfsF0xdyJacboPAwyI7BnaNuBecTOeOK0MhfD8/GZYxGHBb1Ic
5c7MboMaSCvVI1g6HeeoyXMmHQciqO4c6fwhqaYTMLYkQBVsmG+9Ikr92XjrLnog/ivk4QhH2EkO
73/JClgQ1dOjpnjhDH8iKc/khwV7xqETuSVmMgCoRtSbclvRf/5VQPjfdCFYEFhpOu0LORBaeOp+
XIl6U7z3EHKcETfIbSrZKuQXGUxpRNzUM1wzlR93C0qPc6mgRyDDu1REdiAJ/RNopx3k0qICgOzE
e3vYcgoO3KJ8KUw1RaE8lUrWoh0ky3N1rab8qWaL9wfBmyaW40DYERP7OhnbMAvSxoV4b0U64M4c
JxrKnbzbg9AW9TgkUNrzFRvb61vOILrkj0mrdaiS1DWnEX4TP8UAGQmZAbD5bJLB3higWOSrK61e
0hdZhGlcMxl/4Y0V5lLj2/Znjf19z1h0pJIof1HEC6XPTx/+tAWZV37jFkVN7KOzRbpd/NjYe13J
1wwxacIBLrsUOyeky3+QEBwJhTrlF8ijWqwgS09GLF4/+8qMC1Iw9eAwDuZsHD96yUZtN6PngNMe
+1f6OHN3AN28938XnR+A1ZjJcedN5jfCcB0Kuuw70/Y7qxT9Fh5QzXi84IYfjLWGDK9uN0CMIP28
lqAyzknL/GI+kRHf3HhksyMd2eQ+7VEjblanKFRi35xfyWNMQf5lkUNbfaUPGFe342Fk4/+KhIIS
boF4UDUMvxOj0ju3q5Zt1P/MhJ5o1ld3xsMbWpWIvFdc2GsHrJz/seCwvrb90lIcGcTXQWfVEs0J
nv8ksxs/NGCZPuqHUajROrUG/Boa0sFbvz2pMBVEJE2n5kwN3c6UR9x5ahNGMfMQXA03U9bOsLpb
qohiPwfkDAps5w+cQkp9U0p4AI4xstttdnLijlhDfsoiMebkjrJE5TOlNCsDW09WM3e/UrMkTpZv
pcfDs/7i/+ejZZoa/4T6lv93H0DPUy/92imVa2RVDN5OZmHsakX9lt4US5su4X1SYgY+JM5mRRIi
Ar0dRmXoMzzM6PE2B6EdlmXWWtxrhzZEBgwrlzQAqeYtKFQMRHH2hYFsghKb+ee2yCelGQrU90xp
l0li+80TCEe410LB1UDj4amAeAUvBN5AVySE35Wb5cfINgjThS/VIXBCdtGvMxNwKrsfWBbDgvry
QgjKN2Pf7eVXwJ4xTEeFxfThmC42v05DDsEjnAEW1b83E9Fgj5Ye92/YnDx9vcGScHCa/j4s1UTi
AW5oRKDlpvx0syq0GP5vhOI378yUryJFnktvDfV4kUnsGcVb/ZnQN3M5byeJ5lhjKXuvqw9MnNSQ
/VOo2F+XPXjDoEaANQpFeNtd89JVmDgPhh1R3ax0lYuXYrRzQKXqP4Jv0j6505LGTdRQQwosyrLG
clHbGlonqPBtc5NBZFN4Hxd6mMgLkFZ6UgMAxe7mgXGVJlA5s89lafb0weJB0/U1GCHGEKtM5GTA
tIkqUSy5tgntigQ1GZ51Ezem/6sedTZHkZEmyRRxwTuZSgOMNxp/eqY6i5DizwT2h1LKSMmKFHLP
76B4Z/61cfgwnDdXNsdW+gVFcC2ImEr2kRT7VzyK6GtLn59sZ2ueXmDYf/HzknXNH1NydcuSvJ2M
uh4/3Ov2FZCVj0yCNU5YCwuS2wcpEqjrWLP2f7q65zsMe+8awmIFpMaJWht3dSrGv+x1zUi6n+uf
eGX/evB4YngpFGhUdNuydSFHG40lLpQEAYtQpBUJnIADaaoJ45GUB++x++0sDtdVV3uAuDiTwKrp
aQv1c7OxMNquK89ZnLCb6koqwvqqxgqXHoPl4pxst9J9DafM+4nrwxjIeI0iqUkyU9oTrTw6Hjer
wsKaP86YrKZ97H5iRwLch/7Vhys/uqLx0sGsoZvnYL5Y0tyoNi10yA80HwXo6BPNWHBXkMA5hYga
3EKgb0bbFepKtDMqpV9alDTXuNuIcc00q/ZTP/oNMHtc5OSOR2NCWnaLQCBHi3ph4Chr8qbR3phC
Ve8EwuVW3jzY43p+zGAcZlnROX5IJh+nWCDXk97n3Gvjb0IDF9cz2EyGshZMQTRPzQq8TyUiHIYQ
gUbdGBzLKbjxEHvKmcCKKOusze41NEaxooMX6HCDgp0BqfGLT0lH7Pljpqka8MsnVMuQMzv6UoXK
WQIsGR9eLZhYblgJo3kqiKkt9rq/Dr+UvgX6Cf513C2kkEraPVUF2kL+38xWzCrCTlx372FMbfTU
U266GpsXQkKoR/ET+qjo2RpgDXgrxrykKd/OBeoSf6ENMYt0AFPrgf4oQgn7Ey7WA8oNFaXLdvZF
4fL4DFkmsFzgJDxb6v7xmIPw9ZftfLoi5BCC0BlwnoR6z3P8Sw2Tm5YzPThp4vRR6iT9L4ouoEXu
rEAikx04fVO550soKX9rO725y1sFVQs/QicIjHS0WDj+LW+zNdKy0ySNMqkOkusAe2s3sC8Ck1tg
SN4M+RtPGpM25MUgbWaU0Ag8ueELJJ4bZc9pRVZeD02BT9E6OdtAUXKXkd3tLaCe/EtdFNH0Ew3U
Z2Q53KhRzft1r4DIBPcJ92T57hnst4Z9U7ed7XXJbbY7BnrblNiqB+wTMRrdMWR8SmaAIObuNq3/
Wa3hT49Yq/t0Js+0b7dVun2pQSvg8KsMoMTG1EfIEWNKKQk5lQq5sfbqadrQoauN6NyM93HDKXuk
Q/2lFfTYBxFJv+54xtMB91CyXq4mQhFCFtNsyfx0nlj0ZAP8dRJs9g6tNHBMqFX8hVlxujuDSFfP
wFzUR7dpOKtqW8MtLVMOPXQyhPxxXxweRwNHWr/j4owsJYzzn6v3MC7E6TrU2WSsF8ugKL45SxuF
AZaog4k7aJ8++stE+4bQcr/Goe5AHHzTxAjkkmmRGlAYxWGgt29ccBOr1E7AK2FYX8Vf9mm4pao8
qjaxonWOoQu40glH3Ia5YGXc7P6h5LQO08AsfPfJK5NuYCdp6YF0GkPXhDny4Iaq9/VYdVKkw2ma
GQ0PbNJgiiHflPSfs54I7LrsXwP8sgv16zSjbqLNmoeEBBgyEOBhBDXUe6matJNsWu/HVinCJ89l
q0jGdncCMUKoQI6bamkeYo/WJaLbE3TSSTshlW6D5ix8vJyuj1uyuyzQxDTdQUoRHk8h1B/40vB6
tG8eowBq98NOWrIU4ZuI1A0QgZ8l/BXiH8b4Fg/Q50g3BzqJMkSQEdATOhiPT4eEf/TJ0H63ZPmJ
JlEPrCrkKbFrzve2mtdMimGHJQLDbLjSf0EZWhtHukZo3FwlRyEt87jkd9Kb+zVva5aPLgqeKM3X
oopDWKS07AocFd4E49jizc3JCDI+nyXt+yg+D8NMi5Psf6ofvtiqi8YuXHL+F9fBA9fyzl3cGz5P
3DmHzTjKkIXqGbsvkCDFPrBG5BBdYO0dQxIZXzrU1teK9MvT61d6qXX/aRJF9PErl5LUGwfWqk2Y
9ZR3LeMGvL3t6ORIsODA/EUHwy5uUid+ZXtj2z9I+ioeN8kXfspyG39Ac0/NE86d0i4/L31Alo9O
Z+PW/a6JMtZfV0MacKr/TzuG17Jb6ysTkDiB4Q21KXfCA2jfTDiq1WEbsS1s8N0QbGBAjT2dJCwv
TKsuxjnXCzWBCO8g+ZAXlS7IasvagweDKtBIyx2+MhLtG/1lHhBRrmwXWBwnYN0ZAfpyl54Rd7SK
lwwXutU6ReATvC04psxXO5hCxSUHvWocRx66GGuvWqNzen/xKSh2G42eLvaUB4piz6jhIgk5VHIo
R7c1A7MKGl5a+IpR+jOlkh44iqIm9znaJsn75LkWt0xrr+YH9v6li0EolgLQR6xN0cW+CntjqWfv
NTx/bKoXQC5ZWp9raruknS6zlT3HH77Zd4hb1pOZJlTtqdpVpPYwqR8ozEfYw6lH69OsT+1N0MyD
XqM4hx//wguetdzlL3+Xbbar0fiyPbBVuXc7mOSTFuwfeMhLnNq05frtQ8VwjmKevZyENEffoVpI
K4r2mbXGqv9fq7w003Ewmp1Rq/hQUn05m0iDqtmeCiH2a55T7oI2MRsPvfPWjHrP39p1VbuvE0ws
49E84DM/jzNksR/Shisws9isemcyDjCMsGiWZde9ppEYdjXb1wJi1QmNy7hs4vDOdYkCbWAIZK1y
G3t8053FrAJ1/O7cEf5V5oQXd4EtLjE6ze4WPFQkVaD3Tp9uxWr/mmFavWtfn6vvWjT9WrWTrOW7
D7BOeje3LetiJNRwo9zI3n5qB3c7WybM1jdTB2zlYehdOrUThaAraP9qVjwRmWJJy7dGlpqnZ+Ve
Z+6pFupQBPXAYZUZvLqAXrccHAx3fxX9sw2SB0ddZsn621hL1h6eS6sOVEkOb2Z6A5uFqaK2DS3A
oCYb8l4EKq/t8sGlfoEQrlnYSvITIOtTTDxy/KftC27UyM1nFCDakC0tincq4r9fK6jD3/L+fbv6
vBW95f/B7MhiG0aIbEkgRT0tekoooew/ZQqjQFh5W3wdsYVZvrpxOhmzIhL3EqmYth4tJIFpZgNo
SvVRCaJtcLhjZePGkRQ8Oc2jsiWafFR2VPLjUdcJE8xIlJ4jOEdahRnCH3IQvH6D5MqBp3951dtm
iIpQV8XII80X29SkeEeriXPj4B1W9rYRyHNKLh5b6ckymvbk1e4jRbAiDj4Pu3wI1+oFkAiSXG4K
rtvaeEcsnSyEPtpc5Vb5Ep/i9hiuJHeXAAHuUnQXJ48LizKMjY0dQE68R1qOnX+FDZf6fjQuOAYm
3lB3fN4Dw+EX1PE2zZuV+9ZjI+N9n/8nfLs5K8lXKo/hUugV3G3eJiIaBCDjcEu3Y7LCyAfLPsNq
U4piZ7moaOkgkLd4BoeryutGNEhtMq7X3FD2XE+9NAYrs473NhohWgrYnMijzNFNrSWPUg6PSapX
XNnTPSUkC0N48rAekOhhHcVMYnM49ZlwVLHCKhyxdmdsfPSVhiDP3qc25jOtpPso1Nslr3myp/bO
kbJfltZ7eQACUOvlBR4SGtEPLGTxmGQjAIVDvqQjZ6C+dxhDKANaMDNA1QJUEkKnQM93OjXOSkAL
Opy4GVyrnUMgYByZJLmVbnYjMjYImIiXp8RUaEEo8+2u04cWZXBd8TYrMMUHCL/pgU+sMHLR7a4w
tRqztx808EocPvPJtCioCIoUlL1UDpaOJb+8WTaLGPsjztzCc7pS3rr5/0nL/6ZzvuSII+U+oIrO
qQQyggQ+p8ntQi/1Z9LVvyKKyUiTR0AA1LsQ2cJuny+MjpE9Xkyg4ZUbxtsJehFIcK9GnKGimSiN
F9r1cdV3APZJrNM5PIxurS+YVdkPuI2WQmmss8is0Vhf9t3GxGfVo6T5UJ3jfa0hVtmfa6AaDmmq
OMsHbjZ91SWaTt0wOo5NNmzceswT4U8XoqNmblHb/E4Ap50cNKNe+qOYsyUxVJ7axiqWL3Z3JFaV
ermvs1gpTDyEvkAxw8m5O8QSGH158SU8LvHB9n3oPc6AEHTHPvV3Po5pq1x3WrnVx7lHICG3bxSM
pnEES+WhhdiGSdgZDtjqyvz3qwbPljylh/UOo7vR87GYk2d5T8QK2zOHQ3mamlgJ4q8R5IcQOsT+
l5uYq7Liv4RsKbpblcUaEFhj6UKrsMMlT6o7bS81MOpRD2DhW5AmZ30zCLY5XgQhC9o4fYCWt5AT
H1WH6OeCOue9FJV+weSqpnLIeMFn0xa1JuwUy6E2TYN00A33KH6JGPvJ5SVK5FLQRY+0TG1O+ARu
PbjVVr5R2AykZEVGydpm4q6zP/u8p6boEDKI7c2gpz2cuz91fX1IQ3Sysub1fAZupjCm8H/0SZEO
GEByajIpQT+1g0vs3TpQ0Scfw3O8Rp1IJfDENMaZ/X/RGvn9nt8cYbUg/aBLGSwa2qSlSMM6agAW
o4tolrvO0QWLU2fKGnHcP86KTdVPaDirZ5LtdVg5/ztg24TfnFjjhCxGmC6Q95+KfWSdcxWkYYzp
x4T+YkAdPzWVUqZSVBsDuQSZxnJYbvZJcHgdEfsu0owlVZIOasCSFdcuAFPzGQAtkAofzKh8Pmy+
aITbfxbEwARvluuK1PtVK1x57zi2HGckUyTa/IUJRCtjWGCkMNw6CrBgEq8jB1eI6xQB7d9eTtUZ
NX/N82+DswmWzPmGJ1qVLsTZAfG2NIoR8D6TcOgkAqOCAFSrwm1zvNAWQk+HuYEksokFgNuywuI5
gqrxnSpBL+fdt8kzdsiysughJQTGC/SdMazKlU1QJ1zI+7KKWK3tJGEGaqg6Kfjbzl300ZsDBUkH
zZwbgkXRTDPi5AsZKAvMkeMm3QIfCxnZGSrEj83ApQ1zILEHzxngl5TQnWWQYRZHihAQaMoqlgw2
g4lVVp8ILdoqJxHZ7EgLpDw88jEOFTs50CoEgyeuiHsj96tDgy+lvwMtN2/On4uE/wGS44pOYXMp
Jdfr4+Hb/NkhmKKoa19h/8EFGDzrl4IFKlWqROAkQQGLLxJFyqL2mQRkyT4Z9jsIBZCcPysjXs0p
0hWuFuG0iu38X5KnfrayyyiP8droj45fYFDE7rEtfi7kjMUcuGPw5oI+jLEOie+inuzXyjI6r/L4
0EfQmhr9AM60DXCpk514CVt7ItahuTA8k9Es4HCTyh2XAksGycx/Q8yWlzsAsGkOZS8lU+0xBzdU
ko2NNUnumsW6zSqaWTbyqMDQzTaBgqQv9FGDR546Ww6EE7zWG4/+ekO0WpaoEjZZzMad2ffJfagX
ct6d1LcYf4mYx1l1DX9IEZ29z2g+cfneaMR9x+doNibVP5Eka+z/W22+xS3hy8NXTxewIXIepmfc
gdg2b5j/NrRXpeKdXLpR7ikse5dKNvniMFq+/KSGna6B9yG+DqQ2brQI64V4MKZG7OqnSVMvdryB
c+QLuPEfKi7fnX8EKTLGo6EJ6zAmdm5+AVCZ9FfQQyaSQ60IGY8ktNx0UcIeHkjZ1++iTLDp8BIT
dFJsgBGS6FOZ5O7fC+qYj9Mnks/h/bWaFggTH8GJ+b61X6b8HXuYwKGBjA5O25iQmSYO2HpjuyE5
SUkgTodkolAeqtODB/xsjFkNGSxdzb74qICc7vF/qRwy9Rv0dXtnYVf8I3PedNPtKn+/IwI7hOEQ
jbylDUFsAi7B0ZVK4GRLVzobNt9SYxtvng4RdqFOO8730qA7Jz68KkHCeSHfz8D0qSSv6L359u29
6I2ROLygW54Ze2tEoZwnnC7XF4UPdwRs35TsUNwCShsdPFS4jAxPej0vR6haZqkHq6SsTcw0FpBB
JU8VyQKYPTujzixr9GAqqxfL3RdN0djsyHtN/qtCOMI2pBdT3uDLRvR/nyWcWSx2vAdBP/yZIgF2
/z+uQDIQ7EIeJ3+0c9a3OcAhY6Itj/ooggysYOP75a3Rn3LGIQWjO2HcqJ3oX0EdLObauS2f4n+J
Q9PBkdZGt+vwMnMmZA2KMhhkU+8/Xd07N9hbm9XFGvlktEB8uNl0H3GOelDu7pxOkG3JEqjHKKKh
KjloAwl+d2y1hSlEv51XdWtFSYJkbq/QQ5zOi6TnxLMTzNk+YINpylSW7OS2bHXX8bl0UyE1/hg2
faURNOput4y0wDiD3xInnRTs9oIXKxUWwHXNiKE1kSPwUxO1BJsxQ0fZ5jayHa4vk4Oos5096J1B
T++A/20imgldVocV/lVBPH5g4jRiJo7M5nqXItIZuLPlxAo4AAxHcSJyjrygqm35V3fxTWkPSdoC
9bUb0dEqCmRQo84GJZhzHe/nynubhU5OelxSJ/5l8F45IZBl0qPQYGkzuCQ9H1FJ1Mbnbg9OgvAF
FkqhgaBYhmqrSgdWEPzpTXbY00CoF9J4txXVmcD2ynkDCavCCzk0R9eEeTKE8GnRhfOC/kUkj5k2
039QkosxG8XfDftS/7+taMJ+2bhBeZVPW+8tx4eFaHhgY+h4D0wY80SO1s7cN8kZ0gX8fMrKUBsw
+Osvw4PiojwrraAKHhCq+x5omrtN1c8zbKJSA5PPOmFMjZUQQYVIGzUV76+WPzFgrLy5lovWBcmq
XG1QxbBN5EQv7mFeXSKmFeraZ1x5XEhSRDV5Pi6GvETArVh3Ip7Qv5w9Af8jD6dj0qd5l5XgdZsU
X+Nns8EX0TFpoQxnN8DgahHjE2yxX2HwjwIYxTL2qV9qxSJnQjpJftsfsO7QGGU9M9AunO1irVQv
hrjV3DZahCr41tNdZcXVLqbZc+bVT0eb/kIKrN3kM1U/0D4ihRWhbpsY5jSmKDALtNb1w0YmW7xD
72snbfH8mqotKa6FKLoCJMyK3hDEFlTXLH1ggPcW4O2tvL1wen5+u4D6yfL+HoF5cM7n65K3//Kz
SuvTkWVpzI9iB/FlnpHUn23mBRcw0hiZiXhvZO9WP8HwgpARZWLnkkL39SirVK8VsD8X9VC5IILg
1QMa1xLAoXB0ltn37u6JchDWY84EORYVL4wdQ0bfPcv9f4r52lTydmU7RCkK3+ekNxSgItEvPslG
pPzLewMAHls0LVw6aa3IE9Osmlk5N1GW8QpJ6lQmvDsviJenmJrC/ldfqtTXalTjsoBRhYEE6DY0
/mwBLmFwdws7quYRYSaxvQsvI1oPrG/dzlwIosxFswAvQU/dczD30aP2NTKkbdGQGffodtN0nImC
xiIZal4p+WtehAW/BTvYZiVOfnm7ywXs7dCah7WZKGnMu5+7sfSz7/xm9XSIvCOgpGZ9KCa/CKId
7m6+JM4ANv0mtXJQYBMIG0Edwha75jrf6+d8EGxWiOZjr0sTx7tavg5U72FPwAZ//OQMAgdle0mY
neXYsWL7B94G67eF05JEgKP1z/CEg606tldfha+ATCA7Q46KmqiKVWzGRFMWD472+oc8X5NjQZYY
uuFXtph1otxIESRO/FapugowLuxhrd8EK+/ypF8SX7p662pnSdzsfWB233wMeODWrz33TgfI8yFc
bLpN33jCX+5kCdn9RFg6VxhaAO5Mv1Q3YUFGW9RrM4lNJ39xRCF/XtrmDvhY5WFMqh4ya8ZbpFlG
HYaMCoLSdIixDSFzRVqey/s8AqNdNmiMrjXHgVTPFjKwx4roLJbYrDk11fi2AABxyLCDgkdIECle
hvk4Rmy7zhDISVhDhJwXjAxV1gKW3wSpv+GW/vyaJpOaAOGVNhRMhJz8AXzEtIMmEsH5l2fi5l1l
91JhQgAt8IQ/2KM+mE69V8J6D5FgRjaJtCgeSCCJ+mWxzJJ4rPYWadiOwSHSVtMV46STv/xUitGP
XbFN3C9PimGcsV3wps0HooxycuCUtyJvoL19ZKs/5OmMVsgXpsz26v4JBY3TvFVhpJdh04mjDX9Q
jlS724wcH1RuWfbslevFn3NfOnrW/nZNWpvEDIDrVqBeuLjKKW6SCRL3QlxtPaPUH65UNf8wnrU1
41fkpnn2ocHne4kqamnP+az23Y+6h7CuttIhRbR/ivrxQrfeL+KA8webiqdfVrLWDea56W4RgsB6
WFHhmrq18M9+JNyA54NWIsPFBswItsCCG85EyLVcvz2dsJRL46U3ViB7PHSkL4SBtngHZXQ+nHrC
ydDfNc8mrks5ChEhItRPkf2OvYHv9wDdO4j/Xh5ArpIAVCwqazSxFgcRcQeuxFoFDqc53pSqePhT
Hidy17hO7b+vgzKMiwxEJMa6AStNX6t/FqilUOJrI4cRApfXhlPTqzRSBWSZ3JY4iO+QB46PgGHI
TOY0xqSpjY2XSgpJWXd74UnJrp616JkrrRRsMuu65USkhZGsrt7UsCZybX8M1rQOx1xCNZC4/tQg
lKbR0HloGQTZpU1prpsb9jNJqhm5g2slLohxtmzWcLDZUxxw4NHQRTBLghONh1kJK5SJxV+lF287
eJCGg3UlNPG8MgqouPqzigoB/EIEIdfwxpXeiDGkQBYLko+kgb/Ux+/I8bEnKYQizOK78paEpF9/
qyfA4Ao6/eLSPbOHVrM7DBJTJmt3YPbvDiaFvbf5Rz72yQlbpHs1u8W165NWE1RcRpWEs8TMTtbs
jjnaFadrK2JefyrNN1HkdkCPU0NKYSf9h0cR+7ixS1CB4GVJbMOSHndNgRfMUoi+AQDzpwRdYEes
A0BChexRR792Y5HFVMi1LL0WCXFxPHkH8fRMGTDuYtDX0SkJHqhObO6wUzXG4KGVmYp0nnDfqEku
sDwSJOEXp7j6kLBAmzEgrFB5vm4346nr87azjZF3BjiGL3D1My3iDxLRSmgmB90GSXAl8VEXWoXh
9qajofEkLz65czQJ5AruYj/F+0w5Hj0PYaAPRfx/08AVPCoAsMwA+KO78Cn5fUInag88xsyXYtdj
tNHvyU4Kw0wZM9SBTBN3ptzM9+xqIVKezWAcrtOJ4NEmjCzKizfA5yi6bkpqB3Uy/OL1QpoP99dN
l/kikgpx5fhOGo3mwMWqjFugJ4AgaNXzJhjQB6w9RvamEOKvxj642e913tW5h67Z0/kmjiq7BlOl
t9zr4xykVrWBuEvem0UFdCjcLdFoyGuK0pnoktxpSg/1YtEwJ8a/Bof+onY3jZmOc06y2csCwGjW
CGGFA+ZsoUiCHxreAhs6QQPMx9LMLDBg+yUP2Iv54rGDFEF2vsP0Zjw14unPhICNBItMxOpcdYQB
6mb3bOBbiSq8+UD2+B/122D76Ummrik3tIU7cwcFZK8cbEQqwIt2KSMsO0PbVNIgAuxxepb66K3n
cDHviFFyZI4Yj/hhtOu7+XV15LDlVb5ys0L4rs0Qp80hYIftBVpQXNN0C+g5NqjFrrq8w13Om1mP
RyPuz4X1r+tlZM3dP4nRXjsp6Qh4SSaTiUjVahjlATvc148COF7mTz5KZmPOa+9LEN3mQLzFd19r
W7WAzOkERG+0XEoAuKh19XUDagR6+R7Bsz1wibK9ozn83rF4Qh1k0RvOfWr5P6+yBWUuqleKEAhx
A+kGbjFkJsB7fIgvR7mnKus+l5bNckynn/IIQOu2811AR0tiCjouz4TdsCapBRgYHFUqJLdRmHQn
ca3LRrBx2qffV1wgLpkjLPVK/EP72ssT5EdVC79OonFe9Sjr59Qv4aylcEbQcPSKuJRHXDaeAH6a
wtO/SZrNUodTlo6/cakTdl+a54+rgUmWEffqtiQ8C/OyIxhoGyoAwgITCttlhr8OKkils8FbnuXx
bA+tf+VCdWaJ4D27O9hzCT0ZCjcHuvc0z6/3XX5fziyqqU94ZJEHzjTTLL1k7z5V5i+j3vKSZeKA
4d77UXUAm2UGZaHIET84SmYEZmMxYVr5wjxaJYr52GNEOy1soBVfHAGqXgTkelAXIwjesCczTkKN
iGH8+wvop/k6qMS12RzJQ+YD1wSMki0WYrA43OThUs3Z2Jd2iC5nWYr0tw6L+A2YA+rGwVYTPqsf
3nRiscW2KCfajYPJpapz/xYDoWjV5tC+6GuA0wmopCE1pPLwSLlckA3AXrHizVuIonb99NSbykns
srUmsaX76k+SeknaETqZFgLIiDqHP/RSIeCGYYJsk+JOPtUfYJjBlPJOLc+l75ZGddSVPWG3zPgP
XPVJ9Hy54uK8G9ecqgHklT++E7wio+v4F3BWpKyOm9Mpvu/Wh1eqLMwGoyGTf8otIlwjOjf5eLfG
GMr5zzkZUuL8vRltonp3iAiRfdQrF0cHEEKwyhTY1vjyfJNDbpZpHobCu/5nr2Du1gS1VhRtv/vs
2fXlzmo7UbjsG4TwugK1dPcSNr9ST8sZ1t/Ee81CF9zk7Vj5EiC0W5QPr6FG8Y+Hp4OtJgtBLuhA
wkcFI7q2jTBLUrT4NOgQ7PnmZ7/B41Y8Cb/nTIB/y6GPkNeC9DdmNnbhz0XHw4kWwns5ZGDxvm2P
FWcLGsKVOKkMsvciaz2kcQ00DGcxL/xtYOMtTnVbq+rspsetQCx6ysbzJI9hQW9p/t0Ems8Zw9oI
uW/xxjLY8I6UEy05GG6DrUP9YuIqneiQYDBAzZbSw3AIou0GYivA+2NXr7V0rcwu6lCOHlVW6K3m
oU/pu9ZoE8S2HZt2vhjF7GIbu3MW8o2dBkcMw6pdOXptczycJHXOEK52Qf89TzzSwU+lULgB+eBm
uALS0pimtbu71ZkPTFiORkGDNcyPsIKwNZBZ7ruJiCN8+flN66RCn1Txwhez82/xHkUDDAYUVFqL
K0VKBopKQX0owvmx65IoUPTaJlyCKNxAwsELlBxuhYR0t8Qez9eP2I+YDyIK32bpjtmpiXpa66/R
vCpjGWMq+rN8v6Jl/AuA6XdsVpMPpgJkBN+rtmfHGIe7XX8I3QFj+D92nslwV2p0d58WVt0YfbBe
IYL8wEclijhh+Vqfjwour+5rPFeP9xe9AOK1KxvC1/Rj6WCH+LJ4sRK2JvX7E9YHFYTPzX0t9/y/
rMxNpthzKYG7bnnzpycG9hZEX2cVMDA+l6KiY+Y3tyZKsnoLDSY2xLMFX7j5QR0cUC4ZRm5zeigv
Njfs6E5IuUZzez6O6ijrAp93aXUdki6mDuqosysHNEklsr3msldiFm9uS4+v8SbmkPxDtj+HN/jH
Y0Mae+GXMtdQEXbnn6YmS6ryFwxJgmN1hUME0gJYpweXo5yM02sbtiXkldaMeTdrLlZBK9yZzmN5
rkv2CxkCn2zaXddyNoGnLtbs6O1TZuSe0SBZJ/+RY907cm8gqQHWhvKu2DCyEouwWLkrSJXX1bqz
YJ7Kfib/JDdUQ+FXZDOixoyzK9exP3XaCrXzuTgsG+9BbReiAqUxHovcEUWy59O1kHuqEZKoYCaR
oYweu+jZezz8qN15O/8+HBTwvPCHoxM6OeRYtT0DIemJcuZudHjgkQt4rjrPb8QDBw2vbnTSaGVL
jKsjDkrS/SJCaScn1F9mEMDeRpwYFHJ/zVzQzVOzjuF18aQaLYrZKp2joK305eAFu3/eGPyu9p/S
1ehgebCkoWF9s+hlDm49iLQHNQ5GKUbKSX7JeVxLmrOibTxeL1ZDPfM4MpXE+j29PlENJCqZ0kCV
+St0z3hJ5tjDyPTfm++N59so4GzOFuH8T7f1RbqSmPNpsHZkPOYjXUB1JXRavgrLiphpvR3W2zI2
qIXK5Jt8cagjjF9E2Pz8oZgpwfSvReMjSEq4LSzej77qD8+pDcfExeJE0u0t3pWPxbRjqlmMvN5k
4FlN4IyMMCYt9vY9Cff6AQflyFKEuyJmeL78NSCy34lZwaVd44KdYAXPPjhnYfdBNocWv0kBQ9Eg
tv2yfKI+QuC1w901rdfAWEh8b239UzwdWE6Drh4xWgrpoKo4C/9I4aB32zlcekgVW1wyzSbTTmKB
7849LixRkLq/5EeY2EORpudC8VpyCUmevkbmP4ZWbPGucgdI6ut90ZG+H8FvPCOkutvFb39opWdB
8PzuPuXfEboofSTwzy+FAevay2e0INWHmK083U+ymNQrQm094Sp/uIxOtmsStQdqOZCZyYWDb5r2
jEqXoK/laZr7nVQebD3oQ4D/BEFUUj7mos+q02syyVjFcKYijJlsGTc0+AUCXteGV4se/Hqier4p
Y3fEIKrhxq2R3bBBnASHf8XPS2uwZ+4RbiGj5ac9dfq1ayra1PQEPbPHuIqSUDpPytZN6ABsL29H
2fUcRfezgTSKh72YLySYh6JSa4o2PWEILcdb2VjnVCo+OpbtDrs8TB+l+fZEwPWI0DON3PxSIAnz
TwLZQsHlwj8EhC91zTqaALawB+0IzizTfFlVqUVcTBrlgbxl9qUBpYNrMD+2VtrBcbFR4urnn92A
pd4DdW9i8j5TGAyBVaqB66XQ4oFQe8eJHYN/aCwXCv7tfswCaHyehBX7gZa2Py5JDa9Fnl78BTW1
OToeqPbY+MBaFFkYk6bx+NVtwt2iC6jlspahYE7PFtrBRJeOubHy/12MgkCwujOqPPjCzqP5U5xP
PE/zZRZm4vSVCRhFWaDcV4U4epkZ5v+O4Sd1zknzePuNhd2iS0cQjCC8Iz+n74t529nPVRkDm8SH
SSZjiSG5BE9/E5twY68bL6qziRhaMCqjGlfPst9qUEamzgUJJ1+8JJZeGdSkn0ibI+HE9dYSk3ue
r4IOT640nTyisOC6MgC7g0sw9oP6H3ZIvBHNs/gXnsZhLq7cvhOEydGSjiQyQlBV4kOFLEnlOHPa
BgcEsFx7mLxi5X9hwcoKJDATsUlly2NlGOpDIuw07+R/8ZYJeSwf16gycMohYS7XHPH40ktvJVnv
o+yvZ8pL1HgmrY2d1Nskb3uX1i4M50tHmE+uM30eqaLzrVZ8GMAmccAhLGzdBrDW95WgwZpDqWQD
lKUhR9Vdf+xQtPb55x2fCRS02fvwssKhmWF34TLcCCgaGkkqx2W01w1SRZ0zKv86C9h3CHNfn9vi
bEjQfaqeGfCfhTVrqzTuYsmRMqj08NuDjVvFV/4+OfLIgm+r+g2+sa3YAsfrM02z6vp612kOBzsn
t2UfE4GGK5zeBz+c4NaxQyXv4uxsOcjCIYncjjqJP8+8srhEMF69gy59DfISHUvlKxajLNxgiR1k
yJxJvWbgG6jAQVNSXSD51cYgl0af9f2QdQXv4zpTpoflLNeILPnRBm+hHoJAI29RayflwuA7rFyH
WNPwjIRQ1ZNpdWHibayH2mD5Xacs1N4tIVJLOW4K2dBdqd00Lqx7wuWO9YbqaO+Zi8kp7e8EDc/D
DUwYK1OmalNaWcgprGt02a2T6I5ta7sjN48Qw0LsugctVBFPOtC9fXQ2uDDnpPiOQrQVQKwF/GbI
KjhezusFwnVJgIv7aCn1ZrjDo9wEwdfrsvFiVMJauvrp4M+kRH3fard8eIgMA2MNm3XpRZHhutiw
d3ev7TgbwGaqEqgKLAYzo9LwWmzNCXkWps5HTDkBr+x0O+ZT6LbUUbYEuq37Evc25CpcfhvEpUJ/
ztvdRZkVZDlRDiZbzTK7hXbr3+VyzN9rODt+bPDfTtkHHE8aOFJCywWm4i9A5g3XIvxSjP1PIW8m
KxQkCDTv4uZKBgPga0bAM1v+HhY+jGyCT9Be/KuyqltebicOncU8At4pimZAzI2I0B+i1VhvYBu8
wcUrbCvZzcobJVYdp64X04tjyKahEeVni3bMy5hT/8Tcr1DURIYH9oanuViYK5GGignIUTQjQ6CT
T5CLgcK+thSWtH/VB1G9KJysqHhmrzU/f+nDyp/umYm4/dwK9IjPG/dloj5WfJQ/zGIfr/kQGLQs
URNS2DNycMyl/qtN/Ptl0YTYc5AR00wQxcmxWPvn+kR2P56W/VcXbJe3zivGXVRWJ90YQ3obRdzq
VjHzgN0keqD7bYnqarlhgj9z0ZyoYZP3fBjrNN9XNhWbwDXf4mFTGDh3/lyVSg8HNfbVhWZepWrT
Xfr5/4bN2HDnaqsJxyb7+JZ9aazImhWFnp0OgTvVcK8ZeEyQEZN6Yiv8pW4DbhHcNv6J1ZAirZ6/
abVdbI1w4C0MBN/YJjK7S2rxGcCpxPRDzAU42xhDLjer+DqD6Ii0UPtSSi7o4qvUDEi5idMKWAqX
fZUmwR2VGkuwutg3J8Hoofa6uJ+VypGb5qwYm8mpjYSGFso6+lZHDHJp4QlCEF1W6A7VfJmWVoYC
ak/09YL36Oshy8afILLRJ6CteuOVP40BHS2fs3M8CtNzWQxziHtQcz47GG2zh24y07qzdJxoFO4t
u/HQwkRXPSnQ/Asm7ZsJzrThixzoFDruxYsOq+CrEE//mOZ9cv4j9+RLZ9NXPlrZwPJzHlCVr5WV
5WAv6TLd0IFJqn1LHOfC0AMiZ7H5ZOvYi4x7YvPWqr87uGyfpwaPgFqnOd5AdfhbnifO862i2mEh
B9f7jqqKMaV2aruM8ZoRpxzUYvxURgqfby9W1iS7pdJYyrYEugyCEarj6h+AWyRj1qeFZwal9ZHx
ugUdHHEB/xgz5QSYeN399fpSABei/cDMpHnyYmOiGNQvKPuPYMNyr8QoFfwb/JLSBhkGOdgj2iTk
Ido2tYTZwg9R7y8tcKppPhB+uoSekVsV6CO/pHMuUsfM9lstk1WSsWFJ4Rj7UYhCuMPZssAPFu2Z
tNmmRphyqdgHXbW17B9rRwbhpXpwOs84maz8i//nJ9e/ivcggFWsj2EIgZZcjfsqOwTXce7bzEdk
IYPYP7Zr3dkw9UovTsvNLUxuCCDWEkntt/foRg3pNpAksLnT80FReS4jxABvypjNwXSbzo4isLBq
3UsGKTry1pIuPk3tlRQqWh6IdpQqRayolVZwRXoibuAF6T6tXin5ODDrElM3o7CMRUoDgD1/49+P
kWDJVb8B2uv/gakUaYlzqV+9QXqLij7bTQu7yCSwZ6jz8Az1URLaVmBez2PpLtdkbaTHfEEkyIzZ
uvM/RtPsWrPMoP1XDXwtnMvck6fUmx/4QeC7LPCSC4WY6DEHwKEQtTR49cbXSfVuPG3iG4yqhN+C
4HYbPzms7Aad8KM0ku+K1UXobcPkzpueIUUVT4pr1t456q17CFlefW4JzQYlcodXBU3xe2HqOC7L
SkFenA2nWeWAdQQmti6VCLKDfbs382fFHts5fI/twjIdGiOt8KjRUPz74ZA5GP6jQrYytFh1yO3l
hC+nsnTD1zAm1Uhg5oVgd92RQwjiPw6tQdKzBiz001tvC4iC/aKhGpQIDxoQClwllqVF5os4W7T2
j1+J1+CpDmvUhtHXGPNfs9WYO2K3oou524hUni+zdmy0mdjVNqbJGlIGGlAxgVVpLKM+oTcWBlbc
2wHfUfNIrCYGtWoL24B8E2MhLXX4H9Y/CRgOJIhOomraNl4+o+vO3qYj3M8+uj7KLjwRS2w/VmEt
zCj3/fSZWCOmGN+KXsUrwSfVPecUBtKeKNoaOzV8T2ZRBSnXJMNG2I5b4StklOBnFmsmNhF5klUI
pDURw9vKoPFkmVpaEIj+gqGEJR5Yn5nfgLp+KyljedVPtHf1f6sl+aSXyURzsVEPO/wdDqjWzhmP
zz+HPWtwdHePG3pIXehazJBqadRhYBuVCfniR+vbVA/zw58WHdriWV1EX6j7DMZie/NLz9CIw/Gr
yNwm77JUroU7Qg+4hI+j/JVbaxqH3qPnBtflcnSySzuatWXKbetS4rJHApOJXmUDcCArj3CrkBWY
4M4vfec9KzH3Oc43HdUNnj1Z06Zl7ygmSuhwt+oWCh0omiCwt1zXoterplmzbO/dg8Boi6mMOVWW
2L01F3YqHPN2n2X11uLTLkRoCWWihlKEOtYh+8JKYrNIazOXXq0TlG/+3hDUlrvd5ELlgBV4oTQ7
G4v7XeoGoibkeVXLP3Tog3y7kx/MAtHxLuie3ioFyBAvEO9aMyGbMEwydMKLIu0t6gF6L1pzB/J2
QFIQv/2fhO6Dgo0TRxoC72/odrAiS7soi4wmXggPb6D/x5v/DJyYMOga8FBQYeYEUv8gyRP4wy59
PC3yagzYC3mLv/A7/fukV30e1MLV7JngYI3SQBUxmP2dlkj/0M/EkEpF85yo73qTYwoNHDy28A+u
TZqJClZLln4FDxepZXMMrtJy5v0QT5pDioM54hfMG8f9YnG0fxOs57fB221yD6EKecj5eUo61idq
YJ+diHKz7mIBYsiA5yAwOvL/InVl2Ybuytf0a6TEFTDRPeko0RSN2AEd8SF8NPe6NA6mBKtLEgXX
ASUfRIoO3B3DTxjEfZjhxfJ3/+uDM7cFqKJNk8LkzUN9cmI7u+EdhuMKDmSkjp4XLLZT9aA8JPOd
Sej6cu/XCFEyS8FquvxxzudZrlntN0yl9NYwrRGZKq2SOZgTfWNGGnCbnGF+phynPe2dpwf4xPyZ
WFn3BJT7FnM99FKme09Bzjn8PGxHY3a8zBwwz5LspFUZKCSxS/qWoxchvRpV3VP+rQ4w2jkfdNtg
5C0ZE3VCRmY7/3Jic7QVENVuk30Ufw3u+650XimSg3RAKGlckP3Y6+C1GnNBiFCusL2Es+h+vVtN
hUecAc9O4WDT+QRd/aHvXfLAgqx2pyyQraPUhSoA+LYBcMg3GMvPdWcDQ4LkU4Zx16ckiczg0xQc
i8q4nomtelcekHjQIa3YCxFDqSfcIxsZ6xV3TWJMY287FFhT+H1TdxgpRq4k+aSCoCjCPBot7DVn
L6m7SSPgDYmGY7LTKk2YkZPa4Jd3Eac7mRRQ27DDADdhtbP/zoMHMh1G8EtRYI3LX3erGwYJC+ZV
rt7h6Z2ypu1F2uQ2txMtvEQ8g6hhsOPV0UIAyDmzeI2WJR3fAQ48SG2MLl/s3YaczcyH+iey6iCj
c0q6LcWFVpirZUJJVzanUn2Z2a1V0lZD6WU1NcyL0D9eONLROwjQv0JNR9hr77x9HgaJuRnDC1ou
xhMl0q586d0SinnuE2QT8+ebjS5WuCh8/2DIDokWaQJAYtuggkqdVzv+c7rGpWdHgJUyzb/C7gGR
lhvYg2xdfXU51f1tOHhF+X0uj8b8MoDvZSpuZK7DPcyx3O7FizOXnGp4d/1BahkKLxW21i+MU2jW
q3AmBzG4Eudf9/zcCNoSgrZYuriKvegDmuSFvp5Ql1wPZqugWoIwGKBLbXvVocLSJHR4WQre7L4h
+3Ry6Z6IYWWWzekBsF0mk9h8OMV/JjGUMpEVYuCLdGFGBD8grOTdmdkM62tPYoH4PTKGYpTS4bI3
R8a7o8WKC5Uom+7MBbnnnz6+rBK54owJZQaPy7tCHrSoWbjO9bWMjFr7ThnFrFTHWY1KMv1BPsAo
lBRE9SgMOLA2O5t++KlAuO5fF67rUkiLGaqF5EhVxpHUaOMenfSD+GtOVxCsHPPS/GRk2a2M35OP
Er7Fnk3jNgX6JSGyeGqobDG3Q2lP0/GkmDbF6vplDyZ22cixC1dzq6rqo5NwMhZxMh54QSVl3yD+
4LnGW+/Tz66hcxnp6K9ww74JDsL4JxQQqdyV+QJ61DnELawZKSQ1ApyikcQvaIiwYYuN+CgauXUl
cAixZekVoi3+9n3JJDe7RHGHvReZkrZWLUVlf94A9PElabvvzv9RskBwDYzf9uUe1Ge1BEA4dosO
SUeK8fb01V81nb//whXUoMys8dVFRCu750CKNAHt7FkK1MC0HGShchlS2XQxdgcz5jF5f4KKt0qg
gTP4B6joA1juIN7JNwPPnWFLlfXDx5e9ry3M0FJ3lgfLrJ8FfppDJs/3HO6CEp6U2fTtPp95vSA7
5qAdOQ+0bsFf6E/vgx1azo/aGw4rU8/2UlLe+ATgxY+zqOKUYz2LFKVbybCDJhCeuS/ivlWemkui
tuTpma4QvcZN8KsHrmWD0gtwlWSwYWIDBVqO+Zz7s/uJKQ7R6lvNsrTddQchnQAcRFF4FCY4NTGX
jLMrb0D/lYbUK1Adg1y0dZGeYG8iWIqft535tCW9G3R8lWHrlUX1a9O9yY/9VqdeUEyHi/sMF4u3
T4FflX2haIrgKqy/t4TJMrjU0oOWigiLivi32ZWNACAGpwb1tawRdex49SASFxE6g/MIFUFPu21d
YOFd4qNOiXhxuHpOi/qwNTJLPEOw7fAeYiJ5bmEitm0RFwURnGtCH0D2EsK4uGIjxZKaWYuW/EEY
mr1+KWcyNq+jGZp0RQek8eiBWqiVznJ6krNrXB3gyj34uJR73AASxXzg9s5iF4VEy/x1zofheKt5
NvtrPxBQgppIM7e0jjHvJqdEecVwsTt6slfl9nYguPmufZvf82Jpm/3rElpZLWw94sE0Xog4O6mz
tOq0YnC/jEVo3R3c/ceHQeANRmo3/+7lMCF+aDHQzkScA3Nxm4yjg9492lem4zvNEBu3rZkLbBwV
Yd8hXshTZ9rEoVaTw65o1DfPsrv9+wO+fe+PxCpin8Nsvz8mTU07yilqe7/coTKKCmI6OPNufGuA
s9MKQ0jhA/GJVWZKZ5zBgo3u0+r+QP0Xs0dUt0zryPFdIW1G1OaiE8Vt0L+k5BKT1ewOLiY16H1T
HuGkAd8Fs9KvNdBB8t4pUMSpZkh6lKJCZp02f0rWMKkInlHnnUGSI6t/iKLnQ8Q5NaJygiLmpCc8
kbx5yCNj6n+1qWHGeGaTGu4yq8itDVMzH05EBlkgw4wYaLUuHX38/QpPh8bhC99CaaUb5H/SWKYC
FLrTL1o/aS1KaJpxWhzTqHZ/H0Jqna40cX55RN9mEr4i2Ge/Ch9CrKZyayKYny1vRzwNu/zqQfM8
o/EwIxSCYsfcWZjg0YAbjjZtf1JXAyq4fuO8cIoqWrcn9zSVD23qR+JF1sjPTldu+JpFkcW71H+1
bpnY38rq3nXh6hWENex2MC1vi4y+RccDcU3gFJsAT/1AMfSAhpVHq0keZTitKvDtaKHpQdxOY4Gl
j+0dy4rwAKM1p2UNWx6F8RVWdleK1bDfciqQfrsly7ORY5HxfzfMddov8/vsz55cnfVZUsCqyIhy
u9YmCq7gPc+/IXWEf66GS74pcQz/fu2SFqii6jmsk8nyAPE+zyxBgXzJR/6exUAOQohihoWwc8OR
F+ss4XAcDQ/zBTYjWNOrPYHeXnCOKsykPcdsvJPKz0JvSDkplK6jPxRQfndP5qsqUlUEqMX5sRz2
3SZPLmKkAyMsFlThztDf8tQIwdLuL6kSv+Y/2QiGPFxnoIR7fVdFvPTEnVsowY6qtz00JywM26Tm
PbeBCZD/anWK06XxQJTCjstrHeiLCubP6SMGHI0/CF72L8tU0TeiKNw5I18CZmGFPp6dhhhgT3zv
5ScmqFszKFWZCEKupOEhrKmeReOPUOVQM19zQN98TJ2bjrahBGZD4xUb95xslHK4Akq5bU6+Rs73
15WNTcytmmdrkCa/L6byoGNRb6niApQuJ6lBtrDNBcKCaiXjwA/uw/YstSIe99C7GjbX6H3BHTox
8O1ax2hDJTkS9DQGw/bhWpxS6quM18EC1sH4oR/2AGrvnmMh6dVQEiOyH1JQ/SOPoTjGmxGdfbNj
Ezvrq54WgqfcOWSyLzH9veGv5rqP2dMhpatk2rKbk4ULhGuJt+aJcWgbGYjKgT8Tqz3XOnvALLrx
kymFRw5r5mXC+ITj9U7ziK1hEV9tDhO6WVhls05eN4Z6iaP9FLYEepWy4V7NFB7E1j4jCjWtsZIR
NWZtoUPoKELSsHguHQN8gKPNKQzdEUZIvAQUd394LGAZlDaxQYrVsBBvn3EP2J2IFgQI+t+0sDLS
V6evVL+yIKih16E1ZjXJNvnygFY0ghRGn2ODUrGiX9gBI04bb+ONEw3tV7ToFqEpYlCVRvJe8X6E
9ZKgMArYrjp6gaL5p6ThajOVZ6bSPkOncR6CT7U7mJZTtNaVlDLtEi6RXbTTfFLUxW9bof9Y4HCt
jkAOAHQLAVVyKj9qgM3HlWmKOn5hl0B6cF7bMKQzoTun4xGeOjTJY2QDJnkVkfRnyxjH+90xtDC8
4PVqqCbtQ5t2oBgjuB8Fu0SLh11zHCMcf9QSx2CSquyTx7EmenSKPa58kUgHod0E0tuSvyPZ7TuS
DZvpdH78KeUNuN6AlmSnIRb2ILTIeVK6rjwCw1xXFNI2k/wxaLDltTSdLmqevGSBbIXveNvyoBJC
bI1wucRAvoPiktUjIFz1tX2cPcrTTdz+cYtIcuaVJN7MtYp3+KOQ+zKftzFJkC0UGlLVuTw2XmBL
RJJqFPj1ol5gogkNAYAgnKi2vQq6fAGyKCMaL5WPXyTsLDwA7AB0Wo/8BUNC69Buo5GcsW+zPLWm
RMmVFhGsMY5cB6EMLPUZQTMaEPp/1oK0/39p3xnjqMJrVK6L2m6UmbCAB+LEMwHaqzzuMdEYYKV6
1qFW8JrYrH9YHErEbB14Ap/yDffKNUA7AfNqV2yskOfc0/H0RvV3OwGE8VLg8ialSgDSeUlu5/ni
3Hjt0i5OU6X5SMV8nAIOB1AO5wbjlhh3oJOfyG0Hclu64cz4eS7c9PrLMCwcbN9OuxCGJbRdFsq3
hYx+M3EC8N+0wnUQbuXEqqoQ2QMCmkh3KhktGDkV2cBaenMnYIFzc5u5tzsOaWSGNBc68IXmutLE
pC9vJD/y0e4qped3wgAQvcvxx5C5D0M8bej/UbV0d4dijSq2BykHyz5uCOfoE/pRls5ybrMeadoz
83RSMGKqNtJ6qOYZJC4jkOpMTu0LHvMTDhLZK2S6DFfLb7XHk7H2VdO1/rhUeCZ3sfjvyXjKYgd2
4kBKe+rG1oDN0Ot26hsiRRYvkH9IBggM1we9gysGJYPLeb0ZTCChXGyfDXJKt5sR0HyjyIo246zh
TleMa3ly9ItPi58PhHkxoavoEdYgGZovkisiEZyIOCbftjH8Pl+qo7L4vYNguFRPbNRSJ9GnQar/
73TKfeCjjOQn8ohsaZl2xIVqpd51NP22omcNy7Imqb+O+b/PThDyxxJRl4rVKNqizPVUP0HJ5VKh
Rx1o/TwmFtzQZ4uBElmWYu4b3mqJ0Tf6kRTPS/p55LwUU6fNSflOjv0Awiq8yG6cGvqV5q/ILhvh
VOcuK1omMj3HwOgpSc0Ns4UUbxS9pJhh09K2+sM+AjoyLjmEbQ9HjBXOeAmqTt6Czkam+ehhWMp0
QyLuOwFDlf+qrpdLccRfY2YKUZ1KmnvaHMQAu1SgXtRyoTY39OYIBxgVTAf+c8Kqlm6NHGe7LzTR
yyvJivvfWw2DO6pBdtli4QRBvb+jc7jf+NjxC4s4Js2P/Qeybrm1p9xSnR2WKwKbqa3hTPmamo20
NbCn5dzQrdkU6JGq3KJ4ymSpWy2jzWkcs6kN4HwDiFNeS6BQQ0nn6Kn776goNo87VWwU0asi6sEI
adGVPmJVWrsrITQuUJTSk/T/RMXt8zfOjOGFu+Z+aGrkDe8eyUSqcvaKFLfbyGtNeymV4GzVI+Jp
PIeLfV3QoV3F9Ci5xA7e58k92USjTvyUyqa1lWBdhGv9CQM5dBjLJ9RoJJv3WKj4DjEB4t9flLHp
bnTWTB7VyeZkVm9znd4dUHRXaisZ4UCUC5MwfIlfJyE/AtqA5Jl6NcZro2R7QEa2Xm2a6P4RpTrc
4N3GT6XlugR7mVGiYXcBw/g+r7MQ8FRaSobjlbySqOR25atQYgLhOepsOv12Cbj90k6T9mvCtYBD
WH4QbaM3w13skRXUoMe94RIbV4u/+1DRjeW2ftKkVHdUI95gX9CPe1DmPok4bw7UMYOaVD7SsZmi
+2fM9Krwnnoe7UqbZc/pLfT8EAOpbkrjGTRLVqdVPHJ0PPqOu34nfKRtN1CNVPYOWh6TE3c2Qchx
hu9N22QMatl+mV/ThwdfH5EhWm8gcq/52NYgYcwf4YtUXnU+KCQQ0UfEqXbyNi+zYRE/RmgfLdme
GlnxF/FThW56QaPbJnIziyyIRYOIjdQRkVMbKNwKwhD3HasNqn6g0W2xUffLI6oqixy1rlSx+cmM
7T0Of9EtCM7U4ny8qc4AvIfvJXjiv8TS8VuCNppKcvR65hSRDY24CbhpEVGdEwRGfYVmCNXKPYvN
Dr9ksBexn+fjMIEMG+Y+9dt2jGUL7/j+4VIL8hnocT0+dzfqfUH36Bm+BJHKcsMuEUJwT/npHw9f
FBo6FDOu8Vte92jqdxRl4dux53at7MdaGBNX6v5v20NBPoner8Oijfo671fxyxdf3iZkO/X77Tp8
MBIb1dEuK/4HeNv6h1aiv6cZ0hP4V/oemQsVQBUK8827EF/jOz4fgGbXlT6Y4oXYdlK6cTFzDrj7
TLZY/Rizb8bENd+0fCdGRdwyBnsoqx23GwJvI5RBr4w5E4ld3L6YqQZOzIUjBP44aJyBGlxqD4G+
gRra5R3hGEMbEC5jYcStxMFZKi2/+jsDgFY1YgB211sBWZPEDj98wpKyAo2V8UWdYvkyDkq+sPOg
amxBjktSPRm5a2hzHp7+A6iIB1P94Nf+7iuuA4opShCQu9hvntazXpOpeOvvCUsOU7FQC22hQCAp
kjSn2AC6W8pegPAxJqhYZ6tAVyBI0yhtjiAqe9ofVQMuRnRJYYHrUmHT6I+ZGB2F53mG85wAZ+uM
P2nnJFi2DOjZt4tQ4kuBfUCCO0yFzBoxZQ8Br1fHmlFcTesXzvRg+ESjV6+ZCHvIGoJ3eF0UZqmb
AZK4TII+OPNaPLCB9AMSYHZqQEOzTYed1fkviXp0lmquGs0jbKTJ3skhHd7nmbwGVS9ZZ0RpM0bZ
3qjmjRy12SluzC/NwnIf7S49eufLhrEXyt/cAbh+6d8R2WdBivemRX0ZIsDz02NwtAtIOBFeoOb9
GaW50V5rZLuY2J7s2RG6oB+WtUMtzHmNHz5To5aSlGmdOyLkHtjjhXO3UZxwuXN1FUqtIqy9ZuZ9
nKQZ/BxDmaRPU4FGS920mk6Yx5W8OXauu0n2QkA6scDPE0x7HAcFXLkARK5tTbcAQD37XL0dVKoY
280gwtixf7mw+8ILf8s2Ri49IBtVXkRmk1LeTa+R1W1KHYVw8Kf2ACCEiVg1O1xFSbPcsG2xQ8MX
DBODmJ9hA/n6cOBkfHptTh+HSN4IgKTkgs7tFhKLr6zH/Plv5S486hNQiLRalsXiZ7tCRVdw1QNh
xycL1RguInRAcCFgRBHldi57ckkRcmsFONsPZGp2MJcWeYcJVd2H4QUfW0QjcEb0GB3VXdMNzVfM
KogVKrZhtOYMxeQPuNIssXpL0tqMTRJ1/LOb/Fxd14Atp5NFHAqjQCoeVFgQMltNssxR2yWY2AKP
jHAUz9IR/8UFjzXw1ZBR/ZZbPWL0d+C83mlZO9nwK/cKkju3cIwdUOVp9pzKhAcdpf4TV8Zm2Wok
cnQLOUXXYuKxe0CyNb1CWA5zTF7lRcez53k0SD8QjOZYdNA7mEA9SnR0VuSEsevxBfUGpahl/F9/
8ItwPI5e+i8f7ycI6VfnljVIZS+wf7OugkLNauYMEvM7O21lLtRw0j0yTEyiYtnsYdI42MkJwm8Y
LNZTsOdfrmgZZD0aiKMracRLNBhG6Y0PCr6g/8F3zL1IDgB7q7IhrtDYwvlAXepsD6UoUh/pDwkb
+B0lA8UC6L3cvXblTsyXIR2VhI2/9+4DZJI2TnLaUUu80nl3dqW2tusAIOWXwkK6jy7cCeCaQXCq
TenBFOwLEOCsyGzBD2N35s10tqMWzFPCbWz/tdYbbU2JvAYzPMB4U4sntoDSVo0vyyA5y/GgKy/V
R7dghKcCFF0yAlT1ys+9VpQcmXDHwX67YYNLIwrWjEi2EtBPSfssgzWSWEAMUcrgdzofkkdWDnz8
LQLZJ/cfLACqC0dhCxqtd3ZhgW+wiX1ARrDLVxiA8axiqJjN6XvzMzVZtTe5Yg51x2Yffh7L2Q6p
NyjGQpeFzhaQyoChDs22B4kv1RcvX6LcdmHCf04B+yanv+/TPOd7tKZh8d74sqhV6Jkq5h7XAI5J
mrGXG+3kH6vswmKe4px9E/pXdKtr7s7cTslZEqEW6YsDa5hsSj+iTFj/StSlTlSZ9qXJ35NUgc+8
B4hTYGvypSgwb2MEIK5UNS/JZNUr8U7dVZ4XAyKRh8sgJSP5BmOVZvVEfA95Rnp8XKZtPlNiN+fY
+RK75omWKXgoAiRGgDyL5F6lIXxCR8gt4Pn1TA3DDPwS2PQaLPp4uJ6l9vSKROPf4yr51CS1DF3F
H0J/CaXPID9cHxlnTqseMMPjzVgkfJncmS0gWhtrR1jljnq6+AIlnNvID1R+ys25BDUvWHDFEhVe
WnJrN1G5wqDM1iCOU2A79gvimKSchMG14DvRlDcagk2mOIylHbposyGCB1VSNbv0KewWSr6cDmPq
qTgq7WjjZKQFvaZCFha+ATGNmHAyjDJq+eJVkmTooAKPDFMiiOLanpWiFyt+JhyFMgQn8iaV9JXr
pDCN9vOmYICoeFGkucyOkr85ax7ezl7In7IB4tyAOoc8Kwko5vRmROWGlZJ1BBmjK58Y3R4t7Gj5
ZywDwu0uGr0GNKKMX9vHX+w08QHJxgVF+v9MRVtZ6UL0QAbxEELhy1t3ohESwv3pLlY+1/3WbpzG
indD3ASMJsdT4DZJPROu0Q4QtCJz1Q+mVr6R7kkisnlPFvttP5k5+XLbixdyuaEpzeTC6ogTTGAI
xZ4bJrSBTl9gf3/ZnaR4Q7Ly9PY6LMho75QtKVFpNcd6+g+zpXPYrLU5kGp21a/uJi/Rq5Ga1hHi
YlcbWb/WVnROi1zQ9cuLrPhMFqgmpmRqttchqwAISHUlV+78HTr2Lo2YTjPJ9gFAJOgoXWJ0ahi4
rSX9coGsOb3S/HXshSWW1wxEzalqrJ4gRVWWq7CsWAJEW03YFj/zj1Ulv4WiSZDMYMVc28Bv0uZA
MOIl07770iqZe299QXXc19o3tic2ZEtcSjdokZO06CzhXTG758KRvoTGQTFaCUeMdwBgN8RAbe1N
9wtqkmbcwEOZNsg2aRxap95Gfw2sD78DVbg6dzMeTpdQoiK8kr0XuZDxjAYp6wtMrAdv2eDBlH43
RaMOG6yLGTv3VCX8f9UknV3at2qutKsbiQFNK/49uSPEj5QF/TARBKo1cTatqMFa2Q4Z//VyUQdk
/Hig8UMXbtwOdFXDAFc4gViyIJDssGo2PUJwkc2qZ8/obAvyzMOvk5P2mNCJ2A+iBvonBq8lBW8i
Vn/aChGYVtTqt9Fh3jhtlyXByPwc7aNVNhmiDKrGpnqMjL0uG/0hwuL77kJRfP7sQdqi1fdxadRU
e63HNW2vnWmxvCXcOUFpQUsleX9uDr5PrXGpeK8ro2AmmWbhrhlQYJszzJGKGE1rWweLPX1AbZn/
JRnCfsZHx7wUgS9JUlwja52pVMe6nAXqLA+/xs8uWf6mqRKO7OgfCwyAsXxe1LjK1Jmpv3XY9AzK
ieBRfctA9b3mRT+j1k4JCkM8Fv3QUTBAA+yc6F5n7OoEhtD/3Fplk2d2ymOQk0+gdioAKxI12dPq
TPmS7D4Hsmq9W59nPiZRA0wn7yQCqUaWAfKmOk2HUUkrO+yIuIf3uS9oXey9cbZJm6yqX3mMZAEv
2CDRLIeVrcLeGYTNynkFTFCy/W6OUIYa2RKLauKJcWAoLrGLB8Hc9WJd/eSJrQ4SXBZ5cCQ1nEZe
GnOIUo8hS7cLPN6MQ4akbBFjChpFmMqe2BrVm7IN2YPES64oPgJ6/MRqZ1Hnd4IOXXvyBZxUmpYm
XzjYoEvleHOBKXqazRrIAJ+GeZMMCg8AZXdwbeMnY6Hdod9pCzWj8Q9XVWzAOX1BtNfcD3Qk2Bhd
JT6PBAyRCq7mkj+tdLMcwb2FZegUQMt2a/Th/3CD1xwMmF+I2BdDivCvkAJ8ZdEblLGJWaDuik7F
90c97aZAfPqPoAYOzW6T9Aq+A0CG03YbKZjDlIu5zDAN97nrZm/k6KLsREbGb9YehcH/Fsun8Iae
vxnmpv0pcOeN7u2UHgznh0H4M0x5eVRHzv/AGavpXP6i+mRFYZCaDyRpvWaPkDCuRuna5EtHRIWl
nL+GqHolNdf6d0sAnuDDBIBrHGXmx4upRwyXbWohP2XnTvuSAvFYl0xc2zdZnmYzWwY9T6MiWwa2
/zFm6rhG/K3nJqq5nQZUwEw3nZIUBWU8x3ZDHFl2vuRrsUk9xarQ5OIFffK5stS9CYnMOi+l0Wdu
ZJ4W4MNCNd3jWzp7WvivA8OqEaGZ9UhD5bzoN9p+2kdRs6/IOgM1ixIMyKn++qVwvnUeNvUJesqz
fZ5YUzpPunAD0W1cQPf/ZpQ/hvAB198BEAcP6CIar+LREUuy5RXKdH+K2Oe2STu2BgGYPNhWXJtc
RuqB8/eBqOHmuIq+5yPshHyw8I533CJKOskIVN8ephFn30u2R1UB/s3S1XHF78ZOvD03Nyk8+ohW
awGNy5BeHwWiv2Yf5eral1MWjdYM/7XShalcVTH99cykjZA72m4bD5pdOaL+Gl1+7dI9CAaF6J96
WmSAR8oF1ORXVsS+oNHAAX95gYsRnop77gMDZxDRZj/260o/Q+hUUPifgnPbDNhwleCkYnSWB/a0
XiXPY32ndTDhCnE2+6pijqHx2tlhqgiOvU9YSWWUNzbo4J82rkXIl2irSIFgCsGfOZqHY66xO29R
R9i1+f/EgclTmqBAW/MJq+M/lNBEIWgtUqT6N3SDIdMPyB94lc8DSIRxdeT7mNgnpnGxgpQxE2qy
nITNbRKHU3F+V8L4oh/pkVT8wZecYpuEZKTa9IgwabbxShwTqdA/AnqpNmz6M2JatIAJdU98mLwl
ESGb3Vb/vS7B7kAFg8/37JOE8MFAg/gtQbLhKkyn+I3tD8qo42a6obyRbGEYpnvnpLy7lbgT1iJi
l4tYxfLPQoa1j3BKwQKejMt8u9LuXnYDqUSIPrrOnDh3B6eQt5LguL9F9jQMeYXZp/Di2jZv90c6
//xzKdh43XB0DRHPv+mlKWI9b9XCRNmQx1D0e4S8j8dlQK1fSF9douLpBycDghdlpd7V0xYQmOBQ
79ueQ2VfwkAgP2o6bf/VinsSowa4JAr5sEbpKqrUPP5WT/pn81Lw0a81/SnztJKOcvblX3L1qiNG
xHRCBCHMziUF2BCbwJee7HUJS7yaYdcBmNQiq56qrdueloItwJMfRWR0AJIGAZkr2DJlfhE1TZty
q/Xir9ZXiIayxN2j55zF51jLacIcDrHH02qC5UifW2AgSIKXy+McLZwmky6P0tQvwodIthVLz5ZT
bfRVdkePHRIsckW91rBw8CCcIOA8YdT54l7osIj/yyQuG0jEFMdK+u/62eHRZiwk086DNDsrbwQj
p4/uI+1yxJE8Z3lqoLyXQ9Ipx00/9SbEWMpuB6OzD+9ZIO7Blqbu4no8oTkM5vkOjOvZbey6tSKQ
5+qafdYXCYmoGhhB2siLqGwoSmivl3kU5RyIVbcYvm6DOADeii757CjeJ3GT/XZRAMQ0+QsAHAFT
r8Q7zrJi1Jylbm328kPT4jFEwc5Bl28NJP44dYUz4csWRDnSaY7//ILvyGtBjwJ9b8f5X5ckOfBL
aNfoMxzud5ssQ6k58GDA6xP4dkBff9B82BdE0QxtnwoSBZOu26j5QEb6b3llixW/sVfNoaDXyyad
obBphYX4VKIkyxRCzgLjeH2z+oWctxty/MMhlnZ5KoAB7F/fHlnjZBaMeCd1BztzDK4JiPEQm1bq
KUPiKGfgOWw6s64OX7B5NxY0/AqNMeHuOKeoH97uUd8p6G4x5LUxahUHjRDxCF5nIY8mHX7RG1F2
MAwFMLamvH3xBWvTYl4Ca/pUaCwz6jhTbUCeHwQP54Xhh9KIw2fxc+Ik9T65qE+fWqBDIHdp7NXm
Gg0d3NByvgB/yiK9rND9Y7U0SuXbxLsrpNyTS/16EiI2hHVqg4akoJqoddeyZpU1avMMUHHZIovM
HpeG7fEBZ7VI1Tp6n1PigX5p6wzezZV1VR+sxxYCEh8ENgy3ilIKETceoh92zYioSnSGMXoDjTAL
Sx353DhY4yV7XziPO+tIDSz479bwVAvZhLgPpAmGAOKS4JRqdDJFePGnIv8IlNEdHPE8epm1SZKw
Lu7m7ZmAHs1mIO5YQtwVhZL9g8iY4FCbbhdnYKUzcMJosrY+aGZlvUaFGfUmkFkKEFM+/vgQi2AM
24HTvPWQPjqIHoB3Y7s8ybBFwwcLzKS1+wRB1f7Mj+ndTEk4AzLF9M2lU0Y2XVULuzNSjPCh9ICo
4YdE2HpeXqg94P/Xd3hFhoDxEbanNiSbIIvbSru4QBw/6FDwhPy4HF3yK6KE+MCt+QVqkxYPqqSs
9KrEOWdrEU7gSlkU+U3ByhA3fk/1wTsZzvTAT1JjYqG9s4W1XosPdAkUh3La3ieN5nYJzhp4yGEo
hm4jGHm+ip9RE/ZSzkZG9xP35mSK01/cr0BxJQ+7/M1/9RkxEHITbqbvvMyjrOH5z7lZcLDzKqgW
6AnXFtn+AG2tx7KnaBnmuDL0Z55oqzhsLzeZEQTPj/zMWvJ5GSZrSM1m82xfbN5iqgCpGz5r95TO
VxU8QXubPY9gTVJAsdhwUIkQ7iPnTMQnm0pmd1HsxMisDgzRhOVAwmgv5QCgc9hNvTQph68pdEle
Tb6CdATR6a9xSzMe/l/hnY4LkdLpE7kVf78vsMqYYnwlIUiUhXv9it589DjtTzHreyUnr5ynPKCf
2SCMZ5tZkLJ1SYDcvo4f317kZ/LdMTSBvrSX5pIwetSMhD1qbWNElI7ws04WOtaHpgFM9TO9YArj
DFMpbvuNf+9JQGqg7t5ZhK4eBLuuI5g69EZNYX1TFuWM+fLKNxRVPNwmzH+2YnmYH2ZXofbOYp1c
0Yiilx/GvVKJcH1uUdXYvTt2QUNqYM7RpdExk+izoekKjnHDhaZ2Hpyco+XrpF6Gr511akMmH6EQ
yvv4vUnLuYvFhz4nm7Byj4nmd0CxLDbUM6gFzt9LyMSjvUchkLJXWk3Ugojpgo5Zt7Nx7hjXiQyW
eY6dyry3R8BZE/Rj8ixw686g0kc5bvx4rxLP9LRDOGa3jl4JO7CIHmbyTQSNn4MoH07Ax6I20nBi
ggV7e380bytEwxOZL9nVUqAVQe65vxagImEbyP3cwNJ4eQ8uWnr9CkC62X3QiCxfZoqhvc1o4Y2+
3/cSbZDIJBEztvjfE3oDZRC9tIg1TikbhFJ4sU3BzrSgOVk1aeyV2HkunAWnjBmxIaM8OUWrAIxI
iOFL/g+mpa3dnM5HQYcHdVoFdOUEITVyTygYK1bWRFW8UtJYN6kahXzLFXHLcxh+8+CdDfDu+hzS
Ci9MRMus/lL69FTj4Y1L07xxiZWIjosxa3c5IpxhU/M7+cyDQ5cQeeFHUBMwK0qKenPc4cT7RR18
czWhB5rfxN2OstvwtFOWUBa5uH4y2QzLD5Fo7a6aF9aWKyGkiqOcEbSw6XQj5nVa5QBAI7nC362N
aGcgbUbPaj8dxJTTjazI9apElMwtSMrejgGg9cyv+XJ1r6+B0I18VHkMw+5DnunqehCOOyujwg+i
VbF26TOHXyNTyCT36aJKAEEhuv/nX0CBw0m4f+8y6mbJ1MbbPM5wrLz7IZT8l+y4AykiRCgv2kDA
k4+JlNB95ZFut68JUfBUHQttpW/yaynZIPje4uNw5P/JVyJ7ZfF7OQNb1Ji7XUL2y5Wci8Xf5S1f
FKg7Uer2CP9gfZ5pIzi8wfSxwb+nhnyIKFiWDI6ApptM71KG9Yoc24KQTUdbCx5rzz93mS2zmeOO
etoVPrJLXA1/K3WYPyqT9W/nr5JakvMXE2ZacOurwWOsq34iE4oNlcMkBtNqmuNppLruDlnBtuk1
oEuvy3CeSf1pqXzB0oDWMpo9H/UUsdIRO1bTD4AN0pt9PJydFcD9YAJw2DcH57H8DJEH3/71nau0
vN0r7IxtndSEuf8jtww1Ftsp7QCYCPpXI5LT65sysgFr5mWvp3a/+nBEjfq/ioTdSTdbMwJvvJpQ
SYch9f96CtTV15xbVpCSV+/gOogylxhi1Rc8hooNOQ6L/2bIdCqiy8N6Pv3k2ZZOoUgspmJ5Xmnz
lPQ6BgZH/BA9EGQcHofJ7aOIV5Yv37Wc0XXeolJl9V+B2NpKQgvnq6ynPtj8BMT2K6ks2zs9P6qz
UGhhVDXpRsI/63BBzINmcnVAa08l7Pu4MPSOuXF9Ks6y9gHjOzvQRsuMJLY84ITEZBRMP3kiv0/c
Mwa5RB5i8tzGUmPiLSxcgdXfe/JPc/CDJPoM0pZZZXtapAEdm2UwylB/XeTzXhZuKkojf2RSWuKE
NOOdz6bTyAL8GCPF2FlVCiL5mxSRkDSZH1ScqZZ8Zjxx1RzdRXJZ82VCDRWYyOITD57Dlg4n5y7n
8pDM/7eeKWHQeZLm2rydw8dlQtohDkOph9aYbxfpkE9isTCqJkYh6WMNGot/9kxpPCEYk4Zl10Kh
jv6useUZn+RRP12jVHooX33Kh+WPqlFLMWijtMybRpYGCv5hJMcJpBD2WM/Kl6CfMXSCTDRGzbTk
VEeJAP2ffw/RPgRAYv29Qb2l16z3ehfaB1G4KauKFrLYMO6NmDLwy+97eVVdApH4nP26CuzADsuA
PHJ+e2VoZDKB+T93iYzzH7GEfEMryVYu1GbwX3L87ViH366FVg2MirODvM6QjvRq6m4n3CHNMaeP
tqQQIAzded+OHKe1LgJehuVqgCmP70nbjuo37FdhnASNfv+tiCKmZ3dlqi6x7Uc7YkLsSjrICmoW
UTFB93l+kjaxMbX+UjzC8Iq13g3MCpe/Pk1+9PCwLQLBwCsOkppRVGa8Q7uGUcDt/w5tFEuD/ps3
EmQf9O7HAkgNs3h9Gd88j9wpEOC3XHHwPoD3ffPuCh2FA+DjqNPAqFMEEkaLLPcYP6OnINwImMnf
lZJZcamc3WmBu/G8YH+jvMeIHPu66qxhUI3+5blZNp89deZ+ctcZj78Q4/Trm+PfZB98t1MgYvA2
PZm5pkdU+le4pWxVGNjm70VYemWi/dXia5ZnlXYE8lIWYQeljgqMdVaxB8d7nZDN/rFchjPme0cC
pAGZch93myQ540XftG2KJ1VSYyHoeEgRwhn2bhs6vSU4fY3GUWqPfknRJIS4zvhFLPrWVlJWWH2+
bxLONMVqld1MVWWfAEN9k4ITG935MPhW3qrXuAXwo0xM+lQssx8qPpTWUG2glGI5DuKkUFRS2HJW
3yN4UaS2wkLL/MnldpvSQ2r7Xs7DbZEyfnexuzfoLjMZV+DEFMYj1PfxAPfBTuZph5ipuR80Okxa
UdrbezVYTm2vgBftZNsCJXCBeYZKIX3N0XBwOhBBdQMUWj23TYGFdNMz3d78AMx++UMgtbin2uXj
JUD+kkwANLUtVDiFiUl0kHnCEbXsL09CulhDQAiw1Jq4/Gh7ik35yrOqSpDrS3YHdW83gFmYoYDF
XbIi/So22ZuMGUm7LsJSONvd4Ks40PegdDmjPTjIujwfb8eC+1AxjgCbOdQ1oVK/X/nzABk/crWh
HRR7UUFgT1PXR2AA5urXqMKIxWjCA482ThWle+Ezqqw9Z1z2zWMEu0gD7EwfKhoY1WH2c+P1fUdN
/9UC0fdlsUfdZ1PqSin6MqIMrK/eQdBQ0PBLBJ9ApKlIHVJgDm+9MWj19XNqx/3xbrio7FZqvw0P
DbCOA0/cXUzYXWhNFMWBDWaOEafW4cTx4UqPokvlA5Z9mz8OrbxNz6Ng0xGoV+YBfF3ibnBrt224
XVFbMOH91NBdclAjOGRbQoP24Jwf87z4BxLQ8uHB0ITHckZnSskjw0bj0cnUdXnJwQE5OeOdLKQD
ByPV04rQz8aJvzp80x/eg7SGTaQCyzXB52VnHcraqqybUOqH5vfau/nbIGF42dcHzI9QFe/hKAgp
m5mzmydm+H+2VF7Twvdf4dHo1pRjwOxIdmQ7fS/Th3D/GOP9arLjdzpP5yEmuu+TWrb2R0IWj8rG
U6x98BvKolbmeL2yPUd0n3NkNMWto1HiCOseabLK1sKWFyF7LiUFOwqoVZoX/LXB8mYLl4jLpedc
6Y6AaW6YlKFSHre1wMBHNd/Y4VSxTqnudQgAiUF8KOf1IfX6LKFla1Wc8ozRGdNyEjEj1e7XXOJu
8qA0Pb/65VF5/iyqTJIfvRBYQH6W4hB4Gfa0KHc1/zRBJBQatYQy0aNqOMf9eTtHdMgXLF7gVLHq
+cVmby8N+4nLo9FQvVGSSkl16Bd32YtUylfb+LzSdp28HyqoPxTGrIpoM0z+liQcHEYkknqT4Sje
HA6Xh+B8wU0SKLgSuiYVzRj6/KWg1g7Ivgk0zRyHgJUx3KUx+X97ixgLyD+PGfYzYbV+lei4f/FD
ddAFwrUyC97gwSrNAMczxe7BhTgekGTZTLcgFj9ZcKpleNcESkrnjjDoLCaXM8+Fb/c/v0vHZqZ7
kw5zxU2uHATU+RUa+ukEaHQCrq3Ah78Ddzr6GEE0/kyek995djzIf1DwWU2W5JolHWgVrFY0rVeX
KovY+7Ja6aHiAWq1bR2w1ML0hbDXX5Ler9Xwqe4PtwO0tFQpLGkM33STsblYFxQAzl8Wgz7tM2LB
3IO9nPsO2h6Uv6FvxGTjqTeePuMxtqlabqNZ71706+vaL3s03u+KIeaiPPHSRF+lO3gExtNZu2k1
SnLfsL05vLL+sr4adhKLgGnwiDfmw1cF9K/jGYMIdD76bLf58KQDKhKZv+1o1QpQHSasFOgOdjNn
eb0da0hBhUggdFyNNbl5XqK7egZ/nfJUdjZyjoOHcXwgIgDKXOmeZDNYuVOP2Z9fST6uqUhkBknM
LuXMrzgC9aU9QHFlecKVDwiKsJVudsJVfJ9NwRo+L9f5OG87OIerfgCaIyv0D3xIjKGomjHLgG7s
FPqBZce4+PqqX1B0LfXHt1xOP2ZYWx6UPuSPioroTfMOfnO2h6Qcs5UBTnpwFhltrv0E5YXwp/tM
+zlMm/8W8Ew/MAmF3aVCyUS0S91R9pdckXP7/pJbHZgr5FLLq5KzLvUld7EmrunVhCdig15cIGIW
4hMejbPfcRcvynjKuRroJU5sC7kXtYvg20BqExDLphwJI8OTOS3e5pAq7jr+LvdpD1VmxByUSC+C
rd09Wct71WI7ZBEmrYOLPttINSdU0bmgwxwsL8v5iZuBwfcAkUyDk2C2TQ4eels59KhbqFwuOwM5
N2Z9SZhtJQrO9g4q62rERXEhrbxXh5HI2XOXZ6K51NMrh90HuC1qMDI0RB+TB2Z6Es7uE2p2cy+e
JkKtYYf0iSOio5q21g8CryfSzsLofkycSTGAUuPCcevZNQQF+1FowbjJJsFy7j42rjSTVFEEY580
WDhgXERInDvLAc8tt8DQLKkONcIeKF3DpICdd4vqoYslMlO3ZTuG4sYmCzgG3yhVYpiXYRoA7CjQ
EXzHkVKZM6I/es5p7kIFTyi1mpkFv9MmvDaKoPpVgZ5U9sGJCGNe0HR7sBnEwUvOYnxmi5syTO6I
pAdQ7Bx9sXKfjbufRtfBIWBrDPbjKV/z7WKyZvZdTFTIheSHrG8Aa2l6wliB/wJhO/d2fdi9FChY
e+e312Prhv9RYOKWfiLjcJ+dP+A0t4Ctd0eDiSWR/f3aKDOw8RIuSh0R3uKMhsF2KQ5hBxKb5zGD
95QRxw+iAm5zRLzdJ939ilgdAM5QlEBnd5duP9BOAOhQOje4i/LjZsSr6bfJiq3o6QtlSoPFBjOg
5kQkk7yA2y5VTpFBuJ0ytTu4Iqb5AV7xFOcO77dc8AZ2YDDGA4IjOE0rILlXdG1t7fZnxnxA+DIs
CgsaicY2qZC4Q4pKOxW5xPxfkZftPW3iRTXMKfmKdKhRECaA8sQe+cMyBiSrnO17lZ4FLOehyVtn
CPtS5wpkJy55gEjMIPAhkiQu6yTmWHXnSCpkCu40KAsCAVwHWMWaUooRbrYX9VrXxuABi8tPAgMF
77tnyESX8gI23DHW/wp3OrVVFCc4fhNbUJ+t1ZHm7RUPrblUJlTZ2rYa/4vilvjqMWK2liWemxBc
IcAE6Bkr58iwCtgWCqMSY1b6vp8PeNTY4JpTMXVPe9ZKg0/KlNYSQg+ZUUfGS3NuqcC/qCeAZGWG
JceD+sO2GY5+MvAdIJ6cZ0+k54Z2RL0Z5MTFfvaQ5suzPdf6a15v3mTfxgXQajH5cO6sz7d/38gC
hVEezBJE7AQTyLoGFprhK15ofuRU12Uof7yspJSE5lLHHkUELgzACcvmDRmkrkofZFOELUL5pIzD
1BDMAeiUYpIlvlYHUQa142fR5Gdwx09npemEG9S9A9PxwyPzRgNmpXQB8AsB5Wlal3WAMq/9jiR4
RK7rK6+f/QOGznnClrYHyUb6fOPGWIUaBsm6m5HKtG2hxSNfkvmNs7jOETB8WTwKxc04uc/kK3Jt
ffuEDlurB25cHbhUpnKmYcMNBrUcoOFqWVYniI5dApEXupvUDD4t15pX+ufgooXHHDv8mD3RR+8P
o5FVNqBFf5UFchvw7ybTddeVx4FgZDGr6GoG4OhBGBkrazGw29VB5jdaGSa+Pw6K47zX0O3BhyN6
O66UNXwfHsR1ozVdrIiCOkvG+Ik256U0BZtTC9SittETpJGWpYj5mOUoBEDLqTegIpPo02A6hZdV
weRYuztxms+aW97sWwhfsdPgxEwClpxt3Y5HB7NHdebFzaSh0JfLAcmgJp44LdUYWeVcrbHxlYqt
AxYriDePCm+21mygH1YK/Wc1KFmvOsh+I4mfr6uzvGzPPH53JmXdHvAuXN3J/pN/CNJETVo4/3uV
Dlf7fI5RLH0Q0ebMeSU7FAyFWR0U2WZ2NNmFqXO/BI5ewlnQZ3udviwK87zgMOSba7An3GEpAHkK
CTNK+UOGNklxkgE3jSGiUBRDjRHAn5zg6M0nYULQGZ+YRFcS5iAj0ZrXxvUBPEd0P+lR6SV6XlOj
5sx6jTBDaPmyNYJ7v75+fDfKNnXFTRmipfsJN8kBvr+g/ZJlVYA/7xoG+nuqxQ9XO4IF/xTAZ9y0
hj1SyKykRniDV1Mw72tEeXOrNBuYSSNvtwcjRFJj27cPCyjPKfJBEyditoDKEgnfGifWYpz2aPWg
qQ44r2sjxaPXUjyY9vbVKA+mls5rK068gMlwcaxWr4lWhdooXdeqQQkVUtjgFcKhcs6v6JqObH41
6L4zHBfykYsk/8/Il6+jXJZgyy03b4R+/7R53DVqHhugqLLibp3wz3Ud6yNWrbuCZUPB/8ttgQ0e
B1uWuKxT17X+YxgIrPQYN/7sKPhllqmg+ptcKDCC5hNCnpKIsKNXBRa1GbmceZMoIw4SMQUSCPwn
mtACByHmmYenkcPzA/ivcSWOE/iFwJYKAMyURa6fDMEdAUwYMRxWUahBCxsrXexNgDs/xj8piUBL
H4X84qaHy4GpeQmMzJYL+a3jfFZIysjtjLer8qovd0uwNNRp7JHU1OTXT+AXYyWDPAfce87X3T4s
tdatmVOsy6PhrPbIq6BteJZeYUqlpvnGDBtqa0UGtkA4CWoVySHOUTIbviyONc3aRPDJlbp26/gX
+M69NTqIGvAsuFg2Q2U8eyyyG5vD66+gS32xnMPEndAMQC3d80OcTPzp3NfA8R8P/dAiKUGpWD33
T69xTgktzI4mUTrcVbwT3O4KBPo20DqZRI8mrVzleO7Srcxm4+pMQ7hqypKaI5VA3p1Rr8GM3KqO
dD5zxX68AYUbOn694hea613nevx8PRyW989gka9ksTJA6qBGa+lXVWUCTj9A0BDco3nS6xndB28n
wY2vK4Y/LT9b7OWja9K1t46LgD3MZ+4xueRweQ85JDW1Jp2iZ9UjaWIzicpV29E7c7ueZtks9/uW
iXGoaAJZdvEz5KeDOmdxGxTglIvpgVoJhEEiZ0+srVEn7Te9sZQhxvb+tZqjc7GliKA+NSOOb/KG
q5iI8uzTSgg8WSadJBOGbuNaLleT44cpZFdXF+M1hNelO/4WUHeP3/oEJLjJKpGeZ2u6d70bJxbY
U7eQUKuf5YlewMk/H7ZC3pctav8Ap2nlRHNXq2PwxGsZFSVgqqyJMbsID+0BCe3VhmHAkjduCvc4
Xulj5oIav38nReiMKQJnAQM2pKv7oKBgCjzIOAz3xbo6qw+ulfA+lnHSrQQy3LBlKRubR22lxBc6
DRY82cNtZgzbk2uIljBBwT2iqM9mrtz/64lZpl1twcubUE2O9B0aq/y6E7/ITdf1VUah2zprBcDR
cvwgR3K7Dt4YqI7kaCWRY0/rfUQWIUxWqfN9QXFjgQsOVLG1z3EDwljE4Vw4eo972LjVDWca2cJ6
RJTjvriH8j4KwQjT+YQYf36ykthy9FqbUEwQqjbKdJeW1FLwOSWOV/LsL4shB2oki5/EjN01/hJd
r0rprzOeEJqGsR/O4fscwmabofhLAUoRizuOeSCg70/lDoLNcpX6kValY6HgZcZhjkl43Y5KHltB
oiOsqfqDTlnPE3kiqlfKS5Ge6bZhZxSgq8RzoS4gnDtNiV3YZLG7zRSaN4dBlRVzdUeyvjcX/FTb
s/zz0VL2Y7ylolxbCKZzoZyAkKK/JXF0GqK8DQy9L1KTVwODqUvmQY6rYjOFTR3VtqrTq+hPCFaN
wsQL6jXMTvqvWA22sjhiXEPrNGOy7/qDeRJETisNEoEx4vsqEtj0KXyo3zDoHb6pTR0+xIXA9cgN
Nd1KWYp/t6TzACFwBbppFlolw2fUL8JD5YZ//XMvCORlZ/Nhw28NfOw6iwb3Lzgog6Ey1rDNmk9j
hEGYrdAyzVaOqgOMrEe9sebaSz/XHIx5VNzIyChbXbjLDYPTVyQJhLWt/nLYtrorsm72cml4+/ae
KA0gKmyF6OsfDfHU+pzfGFIlb0gCWiBTYZUW2H2lo8tZLHHWdOVZzgDbHL/xf78dHtLGw1EWAHl1
TsOM1QzArDfsur35ulbwL5fO/aWtZlctCgtMUoGZ5Kdo0YHLW76w9WA1IkQtHIXWfBC+1m6HFq5L
qhbVQ+10gRx5iwvxkfrhcXb/gv/64oRGYCDpUXm7OMcAH4WNGM+L5sRaEXV4oPAUem9jvCiqam+9
PlumkFSWjySvlPE//3GaYJqyrris/Ev6UUupEWAM0VYK1MK8Tv9eMtQwh8OMTokBNFvHfUYa43+i
M8ppVWgzE9aO49z6uRZ9Khc2i3GHMvLx7ml/1bIxLGD4TkJJ9XDDup0hz22fbR2FfIKuYgmDrOjd
qW7DnqX6gPQSfGMJTOO0m6dAGRVmlk3CIwrCCRm8zctChrbBDeAOEkNNHdH2K+dUCpMQkkftbKPS
N860r917e6Vp6rn+jIjeIAyK/ZP6eai9LGBwnt0fZttU3yHt/NiESxFIpOG+JmHEPGwkJ4AwZ4yo
967wkdPlVMir7D75qncQhg0h1id5plfRhhVluAxCsAud8FsbR/St24OYnbUwvwWL/fopqo/if7fs
ATnDn/ycJtRcgnu1hJam+Vf5x7hpbVMpcKJsfjoYjaXErSuon6gdtxqs0dTW1g3/XRpRf94H5/e0
kydNNDaKVrc+tOzbqk988EfijnMbS0CRzW/uNXP0QPhjoR3qoYu6BhxVspGFxrQZSud12hcW8+ng
IHxNBdilfeR5nxDFoYlOQMd4Fk9SB7QnvwZVuCNSqpTrWj6u3ZTUxNbMg5mK7dvks7hHhfdt/X0S
04q1LTHzkGEuu+9ikkDxBfjANMdRH4ZcQ37lTj41i4u0DzjX5kmnD03AZjqX6RO9joSe2c6fpF+9
DgIDEAy6iCS7ZcoweKjv0on00vbcxfGL96ZLVdwatCqkfS6BHaCyRH+T6Xryb5UVqI++6PjkrPx2
R8/BPln7cK1YnFX4rkCfIlm6BgVzFJVTggJjtxYEX6Osskv1D4tcS4dA5aDUPyzydgfkIiuz8aA1
3A9JKnr3D4hPTyzp90gBcjiOr06bswkwT4YGocn9P3OShorgQtRtOkf/OJFhxk5M8ZJP1ibujn7t
u4/xoyLIbmIUqrtNsL3R5spsS+EcpzxUQpx310pCKAAFkSAPgWPlqZOkJ2UVU4fPJZu/YqXlBKDz
XVufQaCiRD6eplwufKh8dg1/QR3LyGk3r/KO3yKHqVq6Jvd96CVlKMxliSSR0DIpmqU4vS4HjyQ5
UuUP1oaDp2RtHzcTqBDbxuKNfbalNxdKdINAGsDgU4SLOE7uDHifOLsHfO2xylMIrusQxKpiFKoe
HkRhJ1ZMKQdweWZQCg7wyagVtvSI89L1XGUBY66Wt8JF+xdjpThiJ3KtICOAd2hfT9A0pkIUpgbp
gYJXf/qPA3IkablQexy/Ok72S1sgMLQiToXbMXJLqS2zhqkLEmNTff5gzz1s1q93Gb4zLMkEbB5Z
mz6qz4TauggrExl5p8DNnTtEVV6vw3iNUxKLEukIsfPB9MphWrpfwoxJLEtbSQfMH8VweKxTFf4s
HzrLS2iGcbcZuUwoIL5eLLi8RIRB11EG22GMwpuWiuE1kX1wi81bzcJ5EinBlmJuCM2MZunjH7t3
Ki2gsTiOr9uP2is1pgGSbNIt57ogVcVveaWbZWtNCPsS+mb7T08KquA0G44ZTuRUG6zedZmUHC+B
IQ/t45RCjDDlm8+vVkbwtG41zkuzDKsd2R3MtIqQtF+YWkmeAToq240psvqAndr4mkNJQ5uasDdy
9ckTT1gjaV9f64fLuI9rX8KBa8SMCCLV1h6qFT1MlreKv4AvN363iGIL1TG6U/STacoFljZha4a8
TNJXfoYIB/SeATNddnaipQ2PgUVFjxY/mfpBPUHG6N7hg9lJgFwInXqb8IJCNp2wK/j/RQEROZFO
eFSKq7TTTONXw0zDmGgG5Dz313owm7uCfBEexpLyHvEl/YEdRiREYlRPO183nEF4/O9ZZ3MbLGze
4o0qoS6YBwY79G01FzC1qHAaUMvzQedNpBj2/6txzbQX/+Pp1RdbjUrG4QaRTbQB1pE66v9s/0eO
Kgt/ZtILJsW7VMZbcSrd2npeJuXJ8V59GEYwkJLaBjfG7OrCx4bhd7Em3QZy++wWUkGxC3XLKIRe
L9GYnOITs+Wa+8FOgMdopTjz+oNlHdWaEGzN4+HyStGOiCfBREP70c/PpRYSp+J4OmvCkfbh/5yf
PRYoSYf1dsmGi+LJHbpkhMxrnINKResZOA4eG3cMhz5GbsZRgx+o4Eysd8B8IMcLHQtjnH9p9Q0J
MJ9y0RZ6FPeRimyGndyiOaJrOK58W+zQ4dUD2tfPNVRauNYU/Y1ZXCYqeyHYZ2iSza24PbOBqf7b
7mtAyKhdwlCp5++AZUwzd0QXFMDuw6sAMgXN8yUT/jxDJNA4+WspuWw96THeLyVuYnt7POhrei4D
SRRzICOW5zwkr3mixaqwOgyzIv6Ybd7jtSBCP+DfD/wiMkYrgWhuKLgCrJvrfQbelwKppnxE0zKE
CjIN7b5J7wLYK7kd8mbwdD6Fm2G+rIr5+zBI1kzUE1yxe+4MjBmbx2r0asEZbYs2LSniZMNdb4UJ
XYWSNHXYca6zXaN7wiPVgXE4jQCnBfToNCVvmWf0LTTbG/GP099xseTTi2FSzktBsJthmW7Tv8uH
EHAKOOzzwjOUS9NIqPLbmgnG4/DmMiKK+5uApPtRyxvfnCtFTo8d05Z679y/FtVAu0cr6vrY5ccM
EWKbhNCtMPMBN1zeGgfSChx5cbO3ps6DhOL+1SiD963Yt2jlR+9xf7XS3uWusYFsBIXZBZnFb3at
XthP8AogZX8Fe7YqBciMG9uw1eOfo2MrUmpUrPvvj0jGT8JWTVpNJ8SE3Xpz6uzAatc9axUhxmtX
ylq5OSD3RDxSn/9dVk6JFodakYXXXeL9bjsi9iXAb4ZSSRnI4Tp+Dk3nuOvWUx0xlbTjZ2MSJI+z
0z/bT8yR9jwcBHlT+yd38leGCI7Y7jD+8UrO2UPLN6e6t3YbU7VPjtD5WvwuHbMAuo++G2V0qllk
Cue7SaOgrwLfbeGLEAcNgRuxBvp22eoRTNe+GdJ5DR5vgvLMehCgmKaNaIm80FfmjvyPCFnsVouT
ftCcrArXpwCIO3OOVZY/40Igc7ns159tzSEFqmzFF6QlK0i7sGJISHrLzSV00vfxTo9whdUPUpv5
JGQn8AMYWlPAV/PXH1JHMLWQoZ5ENC6MrMIgqCJWlEWg51Lxwnvw6B5dqAwotjb8m7M/OaRhPZKh
6JYBYUS7yOyjaNiR5QYEgpvX8aRemES4aZqWG+8fORk5dnNSGfpusygsFJWTOEIfm+E2EQ0HEng0
P1n7liIofKJv79s/xlhswwPsPSJ9gLHZgES01hMAoYqvyf5c+F+g8N96LP2sKZKpZIL3d6+EoEhy
M9alUHqwI7Zolj7mRUI/I0ETYstb50A63/lOjh4Hu1KKDJLqBDpfYIPnqX+xl+VTsQU1zKZmLU46
FzJKk8vR3WcyQAAZuYSA+C6t8SjcCyImxk/u4wQWN0i3ZZ/p+dXuA7oaWm7HUqcBFQ6rW+UCRgDw
/vef1ZdqwV8bX96pZ613Hs1RZsjp43PiuDG+5S6d0ovf/NXnQqYkmjNyvQN5Hdrr99ju4J6Yxv2P
HKDZQkMSP5i4B1tZxc0Q7tsCLixYZC9MtQ6YdFD9DAg5SdOM2H6g5r2kKfRHfmE95tjTWzv8j+3S
fWf6QI+YbsnS4gyfB+58eg8NJ+TlHYVYQ9Auu3twuxGlo1awkFXoAvzK5Xt3fhH/bHZ6+gGHh/2p
JBG+Y0sRxmmd7FxLF2Pmci8GxS7b5YCAgsQlQT8ne1s9k2c8EVcgXKnNPSAC/1i4qH9iPYl9RRxC
+WG1YsYtJk1BIKxT46nR/VZ2T2gvsH6cNJsZPfkbPLHyBMQ5g5pE4KragbRh/dQvJMgFl8wjDGi8
e6XrDGmKy6oyQ8Z/5ZqLIktUGQCfPkuZBDJiI4bgjKeY5DXTf7z6h/zYtiQg7ygggM11auxRctB2
zjh4tWfYa+z+NuXpNzM/RIDuY39JbbJ73Lx0pL17z4ga9EsiTqnmg0QxNRzZdOGNFKKdKK4DYpdd
HM1zJoRfnaENcAvByKUGCe5bXScmeyxJbzBObq1+QTqrQ65vDB8vSCC8d6YHfY62mYT2CKyin6LK
laaWgdtaiT8cTtLds1SbgyYJKxutx2vweOEVcLOPNYSOocn4C3MNGLfSyVcbvJMpJrTE8Rk3G10t
W5/eSLl74S/w+fdh7qF6SfPpXHd3OkEy9eZY7LGzyldmbpqf8LSEW//JhcVehbyh7RS8+/FgZjsj
xNz/NRUToKgwjFQ/b9oLB0hEPvH1VSWc3mdDaZSP8uDN538aCXPwU0Y5g5fGwnqwcB0aZZGtRzn3
wjEO73dTCbiYKSbKRxr3dHiK6RpDXNDBqzyHAdpa/3YrF/ObaHekwMUJqMwccFHcMqOv7UzY102Y
dzzsW88Wk+IrDrKrd+uqZM/TTa6wjJDT4gDtQKvoYip4em4pdIyMgf0fgLHazUTn3+u/tmaDUuXa
GExMNeRzQJClpQ2o2IEPgj2Rp/DxhQcbFUuNE0pI0x8V7HiUhpJOEiBYPwJOQKSimGZKilYGzeBM
6D9j1qUzSE2muWNB6j6RNRROq25+cTshHfT0ZCK3xUkh8YujR0wQtyq7Kg3tw+ORSLCU23QF4jGq
YFBVreA1F+19Y2Mdm0JAMLGSqtXkkYfQfFYeFIB1t4omqPhFmpz1gCYyjX5C7+eJp3oQZPAaLI/7
pBS63A0In3FbhCMmvE7ssfMSAi3DvGNnT8K2MGXyAx8wjoR/ni17OLCM9Re1BkplFSAvaCU8O/dq
54MEL6F5k+NlxU/WafS4MeINChcaboi5ZSf5bQomZuOqET7ktbbSChTDDFiFPg3/GVQn0wvYARnH
6irHBhB7VHhgw7hBrXMCFUzuR9P7vh8R7+q8eCyUqprpIPi0zxX89b3yfrQ7Jlr+2PaZcVirxiKc
E9qCvab8reZSRgWGW84O1WsBDDiF85f7p/F4ihFNZWHVBSIyuY2IrYUc8+gPUrpb7Rf7ojsJ+48i
PMce8CxKCgHI914V/CA3TywdJRzBFYuBCnFl4nsoAQpBiHyuY2CrpwmP6dByFOXAAlXj9VuDudeA
q0hqmheM50VZxKARU0BpQgx9yygbuLqAQ21rD0bm4umZzHcJbAXIFWLSFarNl0aCODGp1CTtpfh/
xxAlnBP19aerlgvFMluBADW4GbUka3B5C+Wd7mUyGwDGxTSKcTGmrhNnCFtbfzufZpqN7WiRtVwB
rpWcYku83uxxhzeVxBNuyfi0WM85Yuer9AZTZTgQOTg1Y+Bxp8jOWH7HsMTSpf/YeqEOmFZFpfmR
WFpt3960Ej1TmPVEMcv/A6M1l5v3cGNGel9EPBqZVryOqof+7oQOhtRqQTMdC06Yye0fJPWWQt0Y
N718IqUiJy+ue/x40TTQhMPfGuvmNSTgNT62ft+VYD58vmN/dae/avDW3/Zm/dEEPX32+br4JQ0e
wMtJx+kTSDkaoOvkVf5VP1VSjA7K8PJPL2YiolBV/V43xYs0AXSzu+/Sy67WjCpkoGOcrxp3YPxO
LKPeXd9fnC3rWFQx1uz5dHxCVbEjueHGqPgIQXI9W5NvQxb76CxvlLReu64O0XJfA0WvD5VCe4d6
f+yBFFAzfcwa3IqMAmAAZCcdTPQ2svo8TOSgJYIRveXDCy3qZXTVlhpK1HIOhX+yGbwn+VnFemKK
+A9SHa5VuzdrpAN1vm7xgao0Cxc/RLKjV80rTVNqUU+H8OP8ZUbUS69Jaq2+eSMGGG+c171S/5WP
ZPTvxkXvR02EOIxFLyrS9/PkEZx7tka1mSALFCYN7clDI7vdZhdG05LvyIi2dcNGYnxlM3b4UIl6
5JFn2eMp5bzsEakow2LLKlB4rfbyr2Zah11kaHr0K7VW71pdnXFN0gcvFSptQPONSosEfORDZYGy
vR7Zht8YdpnVbKTWWqsMx30qpX/un+EgfwwNDMFxNDznowbvI6V0p1olRYckJH3pc6rJQ+tkz7ca
G9koAvzUO43yiknRkwDkn5ZYaEfboke16DuWlpMwmq/0Y1rZ8lFu4P3PItlP9K6RjzDGr66rb/yt
O0+y8Ns7kb2DWex8sy/2CqYKXKSdvrPFXHmqnhX4oVAXPr/ZGTY/rhd5VoQOgykQKsXxgZWAnk9I
orGzZece3SmuQEw8Um704alGvme5PrmwTE9yyK82HBZtH6fvQ8GMCmM63yq2C1lJaXAT6pWAL3qH
ocAxL6mFKQsbWvSmMUbCJSYMeG5vD5gt7UoqbTn0nzKR4R4YjGhFYXEU/5mbxxPvOQ7zm2I6Rshr
eHjTI0kM0GHiV5g71yxy+44+6Mcslhy9VUuF7RfNdNB9s3oYo50dcSB36YkponENvnjXclU/o7ds
2kypgsMI3k1l1HJwMK0UwZGS+SjQnF9vCWsCJCRzXjanuFwOFyAs8Dn+J8Rw4SJuSiw0dVMnlxF2
ugBR0NHE1mGRhCKBlywdrj2wB9kkDiZArKHy2DtVxW08+gjY1hQlWjGozBUhopnkMOMdgw9DQhSh
DXeolLz/McLkvMuj26Ty6HCsvXjhC8raKOrx5s0pI8enV98r0WrJ+mcNB+a6+wK+8p3dbj4wuZEs
O39DWmfEBO67x2MHXNF/ncoHobNVzix/28GsvlDbIJVHxVFSVYjhRxaPkRRDAF3l524zE1Atwwat
LjHgsAlB5l5Vxfis9sWD/D1yW9E3WuhxfpmtFC8k3p9sxURl2Z8OTY3RniucQcvdd7xKMofd+K1/
Sw1DDUGpB1kGahjMk22/N2wcIfXno1Ti97E973IGKF7mQMHdbAU1w8kqPpx9nK7gy6ctdALy74GA
Wb+/N8v+X67wGBFyTMqvbbz3gS8H6PiCLZvolkP7OVpknR7viQs+PRoH6lKXR8fTLW47eRAq2D1Q
7z/DSFpGHVL3Ubc5F8eyN/DWOrIwslD32k8MUh3/6Df0LR9buZDZaE0WCJKnV4e8cEkfie8xDure
wJK3HbBEe4VdApW7y7YEjcB6DR+fFX3m2PfCD6NnMxiOPKLjvtyOJALxhr6FmqB16cpLFL7h/Ovt
3aXgQD8tV44A0TLnv3zAXP9jmjsSVgxUN+BXDynh99AwcHrd4JVXkPB2eMVJ6HpzZHddzjrQoyL8
oFj1kiKVLdc3wOfMyjNbwn4HtWf87qo5BvR8YfsOQ5P7/ufhJF+9zMiW8HtRudgoQjB7r6Zc8A2w
WuUkQQ9aIPeO+1dNcuqLLA1eUZEyTjUuRJR0FGSd2oqvrmjqx+LEpVYK2gUHzLtsM5VHwkbiZNDQ
Ky6RdOHUkHYRvxtFSzs7IgE0mygR5vGgukm8ORmxNtiBqo/FTr4zWUVxrrDazjI/jtufAFA/lt8M
y1mLuQaQ+Yvn70KpweBuDDX3pPNMCFpJUR3qCtmwjnir0+23vN13+yU2cd3gGW/tOfc/IPYUCXLt
V/+8qXdJ8qXq6fvBuRvxfLW67XoOHMVTOqeQj07Rs08ZVgASCboTLS3rvws8YS9Lrq8xlaDki/Kb
rdeWazrY+7sT+ZyWRIx5R00Vf/E1rJ1Wt8iUKYF2X9zHmiC34aMWYlIQkJiCCVKIJNxGxMuN521Z
Im4sH2ZUP7IGZVy2dVz8e0Rh6GnoGyOJKNlQaKM+srscreJSbHLtMsFN6d9Bim7xC4tcU7aJ7veQ
ozjbSbVyjl4LYcRK0GOS1HioKBDR1jjTk0ndL/OSyuJCRrgkIfHocMqFq4ETxmX0FrXOYN/hWmOT
yaASkkipr7TbRieJp7dLUhphWdhU+xBshSjHbo2+uhcWCR1WUfAK/H7/gqT/RGEEw1xQ6zw/1EYD
7PhNG1QzDm4TQf41kn7j1ao2cxueRxlqyIT/CEz/63Hq0xQViWZzZ2U+lcW/npvZzO222hc0ybXv
RDBt+chQBw8QNudNX+Wap57VaeuRjKo7RAZGLVVr3GOfpuAN6ETCtq8vZj+JSs8rH9wFCAPWsZUK
rFK+M0kDi/uHmXXQa7gBEuJGMnP7TrmAAP0gKCJO86dWr7GvuRKG6Ylsd6ul7ck8htZCK0LbFDMt
EgoEoD9FHgNwk3adHToRJPhDLx8TBjeG3k/lvnVAEK8CF+5Zuf89h57pXYQj4jhOs1RvIvm3MvAM
B8c3ggw/r3vq9BorivYVIO02e1W33nuDhMIp77l2woY4dhaCNDM8pOxLWHQw69st3CFBp5xrtOUp
8K4lC3R/5h2WKDqJDAcO7WUBT9mto9K2jMxY5bh7iu2ZNZ2YwLihlfCq9blcOgdn8xBaeFEtya/T
0f+ZxQC6ceRUxP0YUfhneVVssFxgaUOek0h8TtQ/u2TpEJRNKvnq9Do+P7qt7l+aUIyUVycL/91k
oQ6MEtiZhguPhfknM/aXeYfTagqqjeeviW4ewahpgzPCcNXLz+J5aqpH2DyB1Tlp/RWyRsH0nzYp
tkEv8Nk3yvL+nLz+on0sW7616fsJfo5SO62X2Sk4jOoJozgk10F+9UdkxAjiLVwxodRX/7qsz9a0
75qTKxYwqdjfzcTWd/8PsUACMKbDUJpUnSVyE//XxXyfpkKRkbHUN2/idvT1ariS2MQ171dJneLC
ugcqTUu2DNSvEE6PMCMmQxPNc+2heUpf0gdOuU17eZzp0iAulMzVhrtTEgsG1DN2ZVkmDmCEi8oO
X79O58WoGXnU6amkuQQbYHuUWmyp91wO66XGNkDSO//itOS9DVp/dnK7Mn0J9uiiZrKjgxksb2dm
UDNBeHilxaRqRAvlAgBT8LrPCANTpLkbvMDXCwfGGrY3HqRCod+B47XGMtus/4KdvQ0exYywAJF3
V1vYfiEzdOFT4fVv7BU7l7Kmbg//MlqmXtZeS88mI9c+FvUZ/RtBVDxc/u4f5BZxtEe+qjP6AAHd
28y6Zt2aQAqS+RYoI1DzgOqx13dPE+qW/obyGh1944nUPdv91ZCIQmZ419RSoT/yrv5mQ5Slm2bZ
VX8VnaLcXZljFvJseVQoPMUjI7nsn9IlKAu/CEX4BAADiPJNIPkRx8PPGwx+BsVzS43CjTK4Qkc3
T4jT7xcj+HAa+6qBP1wajr5RE9i24LTsi+64RL5fEdp3AeOnBL6dHEfpq/Lwl0EZK9QrEOHMxSwP
1SBvh+i7rM0byF1ZzvFqGFseyBxJtHpGO30lQ3rG+PJUkyQ/oi0GIYxTdRrxC5Ah5SFIRKR5tJ+X
ffO2acgSkMxgpO2bSrVyxLD3O58cHtifDdM8ae+7nwwG03HR3X+N4jVsxy6K+cbdUoy4pRwUjpcF
PniJkJmIcXr+NByqy4MeHGiNvOJADCJoeP6PcPVKr7AN6aXyUh9++qXkcckR6MGuuZ2R0pZIj6LB
yfZhTo0d92wQRyF0B7GoDo6ZhpolgzasAC09NJsyRz5spPqEOt7CZbQq2BsUPPpz69CO+P8O1HdP
2dIogzmmiv45wbxvtKdbLUsWzvwjl5OPgWR30xThgd5MGdB3/TjbIFmrTzL8wKdfBnHxuo7dNQ4E
ldCCwsu4t5AtungcPba7iYaEt7SN4psR15R4ujJ6aDaZEMQ+e9ReZf6icMa+O8yGMQnGW83dtlR2
AofmMDgtcUkY8dOLc/JXb/ZQBtylFSIrCqfyt96mlGHY9GhXMPrHSC/GHqQ7qfRjCk04qzBDLWkV
7T0d13htr+5BXNLSTZ7e6rlGoDlcjMqRUBuNFeNhKP+IYwoC7VFxOSxozm9WaawIOIZpAr8QlhKD
S4AicVMVSWtx/LAXAhStCFVFTpVPVSO1s2+1C8Ekw5LoARoR/F04cXMMYifLfMWBmtpNXL0AZ/pU
DkEJE3rwNm6/QtKzmeAdx/72Bl827JewqEKL4rizEe8aofm1IvYuXkQBvcrxsGUPmHgXTkzBaOjH
Ud1eEAaV0RpQUsZkoefcb1LrWKqey3GQO7AJxhtpyjdwvy9SVqfuX/X8hSdtEYzUS3SZe8jtV3rz
1Eewcitk3vc8IUPHHXPYniNd5szw8PLo+fZfZhCHrOEobzeqk8V5+PaSnCtZVqCRN26qVsq/CSxm
n+p8ZZUCKwOUzAJO9yhuo5hFpwkdMlaYlKbfW8jEN9fo4TMm7adtch8gqqXY63Zc6dzjWTBgxFKV
QEaCbaQfZu9URGMTheCadhHxWl3QqGpRVwlPQLX37gLyJ6c8PKXx7gt3hDM6jweeb8NkSFer4ccD
Ugyk2EZz3tLUyqiezND/s7Zm4DV3No8ilRFNQW7Seeo7KlpW92hRh6LBJgI1AItuJKmwCoRLCz5Y
f9L5yE3usgH8E3WHhqoO0dhQPUbcUpl9UciipAWKrdqMvaEz4BLghoVWgT3wsy9CUvzkDb4tPwz4
f6UsBHoHX3bfRtbgha8ZohX7+ySByImLEZjpG4N6rTSIEhRikUsw2C0pavd4NMQyUtZnWNWBD00c
LV/05D1DvLhA3r0LKXSEz86qeXD3jhA9NXgqNrFwC8GcbcAKmU5z/NREF0N1ltArqXfE9kdc3+vT
lTgx6ITEHciuS1S3OEf8lqgO+ZvuiVowXrWdG8CEvqtIgbw6Ok92X5CNvSkDOh45THF0Tod5g+PY
EL5yITy+7AWaD4RWtrNpHY9iloqkmVX1trnuHtsc8+YQSVypIx1MLAQdMsF6ibMLwSNjjMdPCz3Y
IjREOfeu1t+GwVrwFSqshGR17zyvn9RfASJcet8aYfrD1+cekEWZu7tHvGJkQlJSyWzNcccbaUo8
QEo+axUae9FcRWALts0ODA4X+SN/4UwqLJq6eKbu5LbVI5R2gAwCcGJ0QWjaWTWH+HSsV0IujNuz
tLXq+ozEV7KoqTzhfYCyCmgpJO9V4mabw0gqT8P6dj3G+UHRnV8vl+XtpRTViDX2TqVbPKxV6k6v
El8nKo1KBAUuU5tjMXx1tnApoz7xRXku2euLYRjMBwFQqEvUgTI5Ni2j5AZ+uSj3noHkPVGX+HeD
lA3BQohXpTvCuPetWwepM190FyW1ZPSyoJlN6vQa0VY0fCP+9+OBthzdG115nfPLXdgIcHQ5WN4B
kTMuMp1NchAXrHF38blQ7qpjnpBr+zSv/X/84zpbwHJ4uBhOf+XpN3WYsCAt10W7R63LDBIeWavb
/3u4GL5CPeS95ffVhvyKRQ6AmRrKbv+aua6OxBbmyR8nw57DC5RWQfT7Ilg9M4rbUZZmTkiuTm15
5+T4RsdzVPStv78l/dh7Yvc4aviE87PpkzbZsrcWadDuuROzG2yUKFTUFyq22k8GcxyuiejenH9U
yeizGxebc+SFgvkMBxdUIDTQ7i5I9elxNBfF35BmS16OWkj7Hm1o4czoA9ALE0zezW9jTvBKx/BG
rAYnCvKKGIlHnsiaX+C09uzZytP4g6pNB95rXHfE76SXyuAPpacDjPIDMdoe2Zu8cLDoy5lvtmcW
F4Y04CnsY81WhE7VZwcN14CFh+Yt6C/Y07SgqC2sG6PwiGIT3FgBMvsMF+oiSPnHCw+LmgkCveSy
tkyxUcPsNX4CrHQzfq1abis6mvyhDVNQfvfqZYMDkbrssRFESVs6ob8iZCrVU3dAAs/D/6jkUIsP
7HWxy6hnjdmBMKyToEw6Tq253kbw/Um9MJva6L+l5EcMSCk1jHcZ2x1nNWW8hvrBpiNpZFdupwnH
0NKrdg10JS5SRs3H6kVpa9vrJ9aXFs9atjADaB4PX1KBHdLDpQQEaUNN5KZUY2iL1Vmx+nFfT6Jx
F9k+ZaPDWTbEMpQa9n6lGkkBN0CR5Ro957Rx1hfHZFKvI2yDVJLd2rWxEEDI7TZVY9GJ1n+8CTKc
4ie3NpzcHUSF6gJZMU/r7McUrBjAKExbJyqk0kF2/G+qiK3E0rTwsSrrp+FqR8aMNChFVr0sajIH
/vewX7OyrGREyDLNze2YY7zoPYlvI5qUdu1Cwm2/Wxit+dA+CtYDBtguwE1eJUOuMHnWNhq1MBwZ
mnTANRv9on/1/LbkwiInf2PkvcyDr+x2dD9yuoOnjWUBL4fnI1EgEktW3e6wWsfu2hsn81p0APnC
2HZOkX2ZDIYoobfPCrwkwNkU22OWVfpFfSpIPm6AOqfyrZgIfZn/THeCA3ZNkA5Rf/xXA5aDbdtU
2wyrHr2VBEO2+23ximHtqe7M/e6rlksGhHK3RQLqKl8sWBIFCyWaZBKkFg/1rFU7ey92+f//ud7V
JCDD2A98PuxtWVnUeg85WRfvHhCxsLS9ySOXgORVthBwDPKl+OrNcw6MUIjAKNDNQ763blqqkEII
fANou3yuV7pReDmQl70qk9mFD5XydVoHVfHGEtuIDDVNxKSFOXKHOGbQHKxLo4INtLAthPJ91baS
r5IwVbfnpgA2L3Hi5IZCeNixcz9yLsrVCD+RrhUyXkJvkz2kC7IpGI3zG1EA28BxHHCWssXtW7wD
I2JTFiQE0Sa0EWvMzwwv2TUk61F5ABI4LfOcVzjdra2ERH/+LWz6rwsNYQIPc8nI72jDFXgdmQSF
T0IxQSxV2Ukwy7U99NoSDuCd4eYJHXMiO6RTnH+fGR9EyX6e6r317+rsP8jFaKwM2pW3jFFeKn8N
Ug2bfnItgnQaaQOtuXGjJ9hqKoPCdWLk+5v1Emp3YP6u9jsikp1rDXUK6vQdLFwh0pPzrDcbp0aJ
vHxI/sMfTHgfdDOsv4QhcHF//akDKNCXMhmjwZ/duUmtcuHz4wYZZjRZQupAkvB295JkbF0lGCrs
cIYSBoXcj5VDJ0X6YnmTOKSjjCXSmeVOaJddTVOp5TXy3yE+tXIRX1VHV0gUju3EgBHAPx1F8V0m
LdPMrWj6yepZv1RkTAwQyIItW4EOqQ8j/0I18z/hz/Sc2eeO+rUzPOcEPf3YmCuEUjSyZQTHsSwC
usVUSkxWVlv8p8TW36k/4wGdDA20YkadScUK4sZOAk7Nz+bdef6SuHcZacf3IBOQZXKGBEqbb8Wy
qHBqL3IC0UwIDB6d3ZLwzdCIXjsNI2GBtd5WpUVAcaB4pk1mafov6bILoQxGcfuWERK/CmQ9JwTu
hvnpZ4X5bdnBXLx3oTd+eU8fzos6vaaNbZDnzQodV78L3hTJzPrjRgNPS81sKkimvdqDoZF6Y/qE
OU8NlyGd4NNqLg60a6MMyJOvheP8XTBNSgjY4zEK+UZZ7bCR0+FRIuhqsrGMtdaBE6hOoQyeXy0u
Avv3ceCPHoKfPCp/edLzzHn781LrcXoVGrZcBd46aHJZBjmD2YJfR/pd7N+8m9JA4JBbVG4lgUAk
3b+fdDdFcCBlpIUoU6gBoO45Zi3KR72ww7g9l2LU1CJerXfpMc8erxl2anNwOPBq4ConLhG0g0Jx
bfSiYJZVkPjzN5a5jAkEdV8OHMXAOJNBBIQuKkDUOJx7MY0titTNMsoIKQaek9EPq9TRvU3G4yin
yQRJbvzfxnlH4orflS5Tc9sJ8NH+H8COq9L8uBMDvTPXN1+8YdwW82CvVTMMrxLYaxHJgCtGxVpt
DxXTUQko8KPNcbmIUnQ/F+XqtEwivgYV4dcF7LqJU+wwX2tUmGdhGXiqfOwTCCuza1tvOfXl+//E
BdcTFykiEnt3tIJ1lpF28L4GCNiUznWbLnBV9HfGaiQiXaksJC0XDLLB6/sPl+93IW6RAdzaP52X
pd1ZcEQgFerR483oJIH7TAOQPukNeidk9K4pFUlZiz/5otxIJ0T6G40VBKwmgMDAroGxeuLDv4tT
xQ1V+OKidUP5QxteFFrkjbxhZyWVXkNjgNIqvpsBWgsOEgWprmP6QMg/M9CPHvIsnuP9gWi8Zehh
Jx6CYffYpfNqaJkEx5IBbW+O8+oEWPygHHdUq1odlIEtYc8Zw7sxk5UyBxM3rQngE8k1fGzmOlzo
QEvtXfHnnzmLJ2xAasa+/lg2P+cYJ+z6j16i9xf60cNyl1cyMQ4mme+Zu4tmpFSZOsihxmBwDXu/
AqiGKzZVTUlFsEkwAZi63Lqgm1DoiZXUk2ks+q2bgEsDnYoB22LPLxQMTkmksxHqaW4i8fey5QyE
3ej6huWc6LiY3XNaItxtGI1kofW/BG5Aw+OsPzguqv0yYAZA+5XnVOj2g1CbSC0eV0iKTNOtMUPR
z4qgdFCBVDVLmXZuwVU9zrJW13WmarlzplZKDCThtwopMKccwpLWG1uxQdr8QVfZZah09h1PGBZ9
VC480nYZhcEyOm+HmKlzYqxidzwagBnf+N9LZx8uKJsStsc9ogAtH7SJ1Y4gaukdYpUhqjwVwgIN
+U8vqI9qdDq77CeEtOUut65A1BJ9OCrEvOx1oCyhBG1eR8hwlAhhIOWZkZR1eQDfCT+uszqHPqrr
JIBVuMxvKLM3UFj7ZZw+LOadmebAyH+zUN+qZnYdgnu4zflUUdb6M5nQ+g1z0t3GLfFwpt5mWl7x
NvMw1Ab/PM7xAdBKveC0e+MbMNoQZwZUW7qtlLW1L26nTEzsqxq2W9m/CQlG7POgXJF7hLUWo8gt
JD183u2Scx3nEqEsqDpJ2Vgo3bRI6CEntOq4spVJTOWMh44WcIArLNrplnnIEcv3VufbCMiK03iq
9XQ7QwRiu4nEF3u6fArPg9Hvuqy48FfefdT4kVwUoMgUZm2hF6KxoC5xY3Kbmy6GVegQPoSFxB3Z
269mjNpZcZuzZswNo1tUNuzLIL6QXUqIh1CiMOfE5OhCCcPN6+Jw9NO6RM6UiyvDsL6/ZessoJ1Y
bAzP1CkmqM0wfna0m/Rkpc5YMd7rBBMYVfdouMrOpsCnCbbp3EcxawFNPTitaGKUt6qmz7+8YMVO
4gVaOykmI96o68/5zi1oRZ7ZIZvWssAcbGUxzOIsvSAcsL+U87PHu67JdyNSTm0pTJIllJc+7XiR
NvYvW//WmGwA/Ztje8Se3ENIvabIoUtw4aU8jgiOADQDuPh+tC+h52bCjYF4W+T8z7zf2p6CllS9
z5/ah9hV8/WE0zHZdcU7EC4KoSE5qYXwRlulwhkzOqXL98qequ6OrfZcwEPNg7zcZC5R0Ck/jgir
JtzlWTs5GNK4fHcmnB9IeHiXyqF00kdPvYV+WxsmVAeMAI3g7yzhDTCTRXvH8AfPPyP2tiWCZgQD
gQoH5hknRf/TyP+xMz/iCF26CGFLHcGrO1hGGGqjm9CyhJJ/O5P5E3A2J9EwQUhAZPda8xOH94iO
eHNBXuXP23xJNndmQb2nwqmWlZxDh8MI8KynlSJ/aQkNNTQfJBJEgXarkxvG+peqx6M9skSaPwye
gox68smljHNQCU9Jr2eRQ4RzbBTYXi5G/DGDpk4xM3IOMiYQpJK5S3gR6TIZnHwXO/O6dV4YNCKw
Hfx6Z4pQYB3wkKahNsoyB2uBLmkiJki0kFKDK+7tIKUXtuu4mqaMA7oRTPmr8oe50et/A+crSOhM
StLQQuYzGAruCxrVbYSjQjEKXF/Rcegnk8JF38pDYJFOgqz3sCqSp93IpqWtM8CGm1ADE3L1yEcZ
Sxj5wfJUovSo8eW38aChsta/Ie2o98GGobAfoH+P8xG5Ejjv0t038wkASUv+cIr+eI0sZXO+XuFz
zav005nnWYfJn/Zc6jATS8T62QYkgP2ylvd0KAZOtbHuXZtyZwOVFVkqv+CdJv9jUoZMRgR19Qwo
GB3SeW++cR09nm5tw2KX5TIvQ4z7KVj4HOuG3LCV/qVum6If4XWWtIneM+RuNJYwSFied0ZIcnKY
J154V6lAQyOD58B1Ray2rxHG6/CEkHd/FkB4la186nAQ0NOqzpHqW9CxaCbWNpfeqNgzNOSqQxcN
OfU6DiourbCuXdbMPpsoHm1Vh4HeLgrHZjmwpdghFlI/JAf9f2GDJbDAozex2mgLdbPlObeUDY0K
Rd0qlBXOnQ93T5aUIdnu8fYQ5Vbu8mMgWknUg1PzJ8si0cUo84emQW6/Z0hiwZ0V/cGZeLYLJPDw
VCXk6P7RkxQAh++EcdL2/UTjKSMv1y8m+2yXNRkdYZ8iccdV4FkJKU16f+Nkjfek3JYaS9XPp5Yf
raV8EQXKuH95/UrD60tHqEEVKCyMqDkOMw7Y0lehlquzkzGvHvVBlYMazGBZ8I3Vh1Yh+dyYRLxk
+ml6sVpO7PcfjYwbAfGaWt8e3iZprfp5MZy0IATo2FFHsdLqvVye2DwSTDvXN4SLq0EWcuVA4f1G
kslcwy1gJmuaeFahiyw0tmybl9WU+rem5t4hkZBsouZL0Jo1eQ4Ztz74iidZdexV3qHwQIaNSXe4
Ane9Y1DMEDOB0R1VwRMsxY89eH00D9e0tNxB2Nf4peNB9CJ7nKxl/I6U/0+Dcjw7pQxdkkCl9JWk
FM4KC1XjQn6mtX0a9Y7wNHSOh0T6+ksuhNiQCOce1xysz/kDPn/Svi7VdSNSOLbVfqXbmbv7RPWE
/8SFS4gtW43QbLTdI4TfOJrUGZ3h6ZFx68fUoV8RaerOejzxTAT6FanZW0l8fm9gVAndQECaO2LI
5X7gAMJIaPgTf1MLHoabz4o8YqcfOdjmNjnZR6L09NpAj/oUDhiTR9KwB9fltFnpdmFlOBVsac1K
kGJ4QJhF9z+vnAlzwIUWM+vr4w6e+Zhyp4yHyYfolAm9IOFPGbhYhPxKw5kP+rdg2Dnud8egHmGk
zNMKOGkBtDf4tr1S3hhJrPmTiPuLu8UXRZh5/08tyXbtDpViek3OSHViEv8YUWAw0HiuKegKJ6xb
TqJrPLEJ2qZHAMQNmOZ4lOPhx8QbSEx57iNdCjoNb3xGhWHpRK77tGEjKFDqcJ2K4v1vTgTapvcs
QnpvDV6PeG/ev8jYh7JnbCTBocbWtLuivmrvCMFBG4XYW7ye6ij74Nj1dalmH6IFDij/FGL79Ltv
64TMpyYxemjzSqRHCW6zpCvkxctK8ECJMkkPfyMd61tSmX3Y+3ytFS3NmUPK0XBPAAGhlKxMt7bQ
V/G6cBCTMsxMSK3sDW62QDnnDGZgPW7+mj8pSOB23SMXFidvrW2TPBLkXcinqgBOrnZ0UZBebrtb
Fb6uzsXSByBgwNtTRR10ZhozHXjaEd6FOC0pIJRVJzlCePnDtfgsKFHgdKzw9MLr/J35Xk2VfLka
UZQ8IvJi703MGDdy+eHYtWfPiAC61jV7SP31E4vvljtLmtQEJ7NamBalq4WF7FPudfSnAeUKyLlR
edBEZdMqK+7cv+CSOT+ywYyE6y+W7MB5m7xZS3WpnnM78seVOZ7VIcnCNk81Q3n5Ut5Do4fmkGww
KCVDPOAGhrHP+k9CNEpOP5/9rpwW9hj9HziEXh8Vvz9FsPFet327lqouD+IPANyC+K2IjM3mBkEc
U3UyS0oiGyVdrcnuEABIUTAXiX1bTUeYRwyIzfU3CKXfPuiQ5xbMCDQVREoDa6huIssigjngZARw
86OetjTPudHgW2UAxDQUA0hVcEPYvdfBwZCwbyK5w4y4vH6eiGBy0MWLqqXeyt6lnvAmRTigv0AU
GihAuo/yVLLzCFaE4VjUBzlBnY/boPnhK4jqCox2OlKlmIFrc5B5Nnkj3GHVx5Hcx66qiT3eNEjd
K3WPr6D+61pkzjfK2lhvN7T13YYeLCrxJGZFNxv1VrerNI4NOPug3dgQw0iQksMW3/vM2HkqBJMF
J2gTb2o01GohEv5a9a8ULw1HAEmdBBaefzUWC21eAYvyhMVuP+egy4+SnRLecpVTy8K6xt/UdMM3
9ZZdoIQpXrngyG9znmprIzTHEnN38k/pUSIqDrlm48jagP90cdsWSQ+Z9SB3O5TMK5QyjoKjIjXw
Ljv3VcFzt9SOXTHUWg3rSSG1IF+7jcPZ7Zi4uRB86olU/Se8YjVElvSg9rC8B98zepcIvTtVsRPu
kv1fQTs9/tGYNeUzRzE7V+wBgsWP3Zlg/G1gRYSl7/DlNwHU228yMiTx0LwEHPdsyRNITYRVD78m
xVwun90r8REehXj6cNmKE1TKjYCguRTQzSojyqSZResooJWlbNlPwFevMd3FjepW8Mwiw5HdyAzQ
ih3Z7x2ROm14knOglYueGfjvyCPZ21O4SA8AQm1r9Yb/u+5cHdn7w2L1VpkHnz3zKjKazm1mTWAW
thJLSlfCqLNPUxj0cm7MigWJM0POl2blt13F61PovW7JBaxW5u3bgmjH1cGPVE/qMUL3V3p43vU5
q6qwtCTjUORkZixd8L2Ui4nMEOUHjiVrxnqx+AlCbi+e4CfhXMPva16VBs6AfM0zDcXpgVTZiu1P
LrGok8a7fa0044A47zzF0pC9K/WNUFFH1xUQenTcZzZB6SaZTax7hY17PBHgKkKG/lXQYZ52ebYa
kuO5lQY8PikMktTH3m7iAY6afbofGLdCXQy3Ykz/ICMuICH0e4KqT4nqh9U5zviqdkeFKRGNvQ0+
LHw9jKWBy/OPxzCaezJ5uIptpMTD7cJm44NDXpHKcVp7NFCQ84/F5KMCN1zveNP4mLnFcdkw+MAQ
owok6bb837D8UMJE2I94aqg6mB+opC+V7oww+mYWyl/OIk9gYD+x+Mz/7BK2vg7/Km8XY9kAEPEt
eqRwgA9Xwos4jtwOdJwVzb2y9N+7fWIRmo0UQTF96UeaE5Nlv4eHTEdADJe6uXNF/24UYquI1o8P
bLG6FxS3/2xi7BbVZyKxz7KW2gNK2zkpNG7aGpRZu1i4DdxzdJ1gBL3T6d4+uA3XpY/nkz9eWE9l
D/7JlxmNL6cTni1GiqfoMGpD7sKc0ETnrAVUe2AIRU1xDUdTEHwcq9yIocxLXgfwdPwhkKIfe/QV
aWWAjh8imWRL47BEcwRARpFl0731RqhvfZrB931rkGI6p1C0D/awJyQoaIfVpAWWdSzWQGnqrdN0
+ynXfRcAmlnef2RSGwVDxjAz/u7T2Nh9DwGlhtIEst6CAoKeopc6VSOub6k65DWkaaCNxeQfjzXL
CV+vPR2voOOLPO/o93ZGuTdZvhZ6y8iEEScir4XWRcafn3hNNuXuP+rTGq9zh3GX3HcBNiPvbWOL
vVkJFzupVOWFQRiUc/40eQS+22aTU96oBleFAEStCvbs1nH8sEelHmzF4fPsTNJhQjU6kTDyjXzd
6FZHcC+giQvKwjYF8gZVAJdS/vRPUvBPhW8V2G8MZsW6X7K2qg3OFSxAnARxnvvfGnT70+g+oVag
WVwuxpSQFSKwATBd9eoRqYwHjxfD5DRop+pxZ+rFeR7u2xBQEARdKNB9d/fVAQnEZr6ltntW7hQa
SFsDq/cq5XzpNz79e3cJQUjhDslVgC9BDXBCqOvheZOjS5dDb2UukBuU5/akXqZgL0rvxVH1Guc6
KdZ+Se/gnbXFL91v/8Xl3t5jP74cglFIz8SnFDeJpbgxnaf11lsxehB2SYm3LVdjK+1xUTouqNEf
dbsIRlsBVBKcmx8rh2kPAqp4aFyodL3ZOb0OkMh6DopIXHCxChcF+spxqLf5FTEklzza8/4EPFLq
gNGjxDynKQi2LI0Q5fU5hh1nZe8Xc/8+Hg+QSAvNrgDeR/ZHcH5l6cOTvQbdS4leCOoYipRZKbSs
osWhlh5oxhSr7/3wfu3EQA05Leg+K9Sn6kpeMNagsgFPfQj6TX0PNYC18l+OsuPpB7e4mDGqObrB
EavnpQXFCqKh868BO/458AcU/8HyUsBaqLJRdtnyK3w9mjZlWos1fTTM3Fvzgy1Ur8oxx99D3iWs
sdH7kIzERQoRTINOCKVdv49PDUJNj1lfvrFVzv2IiaKVkZYYqy/6W9RluHeVAfsWxhkTD+n816+R
5LZ2Bs8rhgxoHJSIOVeua95VHX0ifeJBX0dkZAdmjfjuTbfFxruUsl+AAgwkhICAtpetnN2rCxmy
i+6ZMisYHIOvYkVIXfttkFfjqLdiQlhc7zHsB5CXG3XCsAjlUYZoDgZ90ujTreproD8pq93C48FK
k4Q/0ec+Uj1vnASiqde8AfY/FKs+zRUJrHr03ZRUlDx0jni33WUKx3hfg243y9a1mqd4aIAGBv7o
Hyid1AYeagY0ABWaDMN8zvwlOm2Q4dqEpoX9rHxnj+R4miXE+TCEzotP6UrAW6XN3h/TEholLj/2
NTXOeOpCCIuastZgIxS1IE9SuPTVy55jwif5nDHEMVeNdk3cWd/QbEGykKfPYX90D4gojT8BIap+
FWeGVZey7yS4gMXwG932K0pVT+xZ+iifalD7Ax3FVwxUxAVFK57W1Ox0AW7Wk2EoZi303KWTsYNk
M1BHEA9btQXfym9NBbFHaRgq8b8nuwRYCQBl7g/QZ8bulN9iwrxd4eZmyE5BJ3zxtkxzco7pEl4h
Wm/Zvf15aN+/GNQ9prtiovBUzaabh1xFdQJ7c943KT30vQOzjXWLrWkdDf1/4724vh8ZTc7DELuI
QMQw6xk0L5Gl1l2xmtshEQJ0xzkV33H+L51nG+tUTt8PvSCGcE39HOEls0B2Bw/e+3mIOq3TM/zH
m3S++WIEqUfWggLiR8kcm6cZGFaNh73NUoyilPmMWG5BvK7hLYvTEUx6o6fTb9iVighHYGBXCj1N
xJFdRKJw+B5vUPYJp9Fgzm7zZ3RQ2gzrRCnZ9rW2TVQCBQaDBI+8KHQy/Ogarc5m+2BwaJN8kEkZ
tPcq3QafUhp6elw2oDcRBjTtNLZgLKYyg0cUi6/wI7YjUqq4sGHeJFnpL93p00BEvWzZfZ5DVXXM
ACjGGxAMUGPyElX0tN5b43JVoAHCkluR6+DXEHklCSeUc5yodtwCiCLbjoLr24EWWX8fFUZBcfJv
qfS3Mv54ZJjX1oGsxHQEJO8k8FV8xraD10kU9qyWLMGTtbBxK10cXbzZCrAU3PvCoGPzmovhiIus
BAUBfvPdjFSGQLmZ+gz4siYAB5WqdFrNfE5POQS0Y1wJAELlt7Vp4FVZQW9boC4+dgYeH7cmQZ4b
79JphjaXZBXIobHVFEaUsE94RX8dZv/a2c1rAwFxhd/e4pPBlYwZphr+gQ2UaFK2yXVZ5IF4Y2D3
/8nbY8uCuCK71moBLAf9CT0lRyC8qsDloy8sA+JLz2l4ecW94RgaljEi71Rhy80kW2YpR8LzYvRJ
+gNU7l4+Vqy6nliHs6pC0YyU9zQHzNwH4OI1ABfn34dcUVxIsUTwVkmbmE1xRErYeGPujbwL1AQx
3zaPwq5gtrOj6rkYDKMFCfsPYRlURsv8xnAr+LLq3RBiJ9QdFMhkaL0qFdRzpPlrV2rJeQ/7nKel
boWoOnt8+UcjDf+VGGQGBraYHvZefR4nLynHVSIFd2PAPBwIriT9Wdab4BofjNwZvRHCLqX+LsLl
BrKb0mTheOKw2A3GZal/dgkTtMcA5jQaWa8pXrQ6LFIjw5n5QLFf1kglAw/B0MykAilK5/hjUBbM
sIX+94OdERufZ/LfLGKpb9iIobNPf+2NrVD62eGwB5PW8M5IqBnes7YZnKOTB0OOSB84hyewD2WB
aahOLDvsW2zaa5Sbp/sRZgYlVPmkYyJsk8uqhB4h/Nbgcy+5UYiz0W+lVfmddyoX3WUFgH6wA929
DDSrarXR3xnlNsIaTCO/oTN29WwtzxM13CZXbFLU70e59lVguurzS/Rb41+JMhDNshyZ4/oe1ByH
cyuSa255rWV+lEkUi2StYL5L8SHxNOAZxPn4+9ad2Ahv2mv8PCffKd5PLYB8HaARAGZimcs13lbR
9GfhJx6pAfgcJWyXsnL8ws0NozG7lxiZhhJ0Qdszap/2U3O8u8QXeid3ohBSsVfcv9/FvBrgFNCR
NwJnrMsiLHbOj2GRaah5Ahz3/FUv7b1/MyaqFmQbeyzhJcw58EwFoUBzYBFFDHAWbaxjtMcGf17c
QdEEvExHTRDkwk9Io2MvqAA6jTyzbLQcajoguFbMyTfdkQuihBFVYUGk65Z8HOIAJGiOmHdiGwiv
L2C/jTUT8UJKXqflRMRnbmaVUvwpA0I+NdkVHFDs0SsspT/H9cPmp2/utmp3fXEmHYJ1pR5yVO8B
G4G8/4WBFnQpctWEs7zEw0v0Yh7jW2ZXyyCKfdyiACfyrDo8gNEwJykIbIgXo84lG79mUYjrfMcc
gN2W6rct4W9xiXQPCk7X1yQdNVGZVlK7ZrsafwP/f5fuSz1/52LNhOK3ZVo/jkLc98K3+38tTBqa
xS4FQh3winmUYRFkfvrN/NP9zTQuQIzzqSeSHXsO1JC2ivLTkQ7fRRgCwtw/YalroOExaYcIqls8
Ucba+GAQ9lAK8YFFCN+yj/euNJ8iyGUHty5pL5QtAIhocBf/f9VWPGGwwvDncpeFyxtg48j6pejG
rGleL60yxXjMauFC2XCibh/ilb1UZrKAqR4Ml2k+Fc6fYbpnvCCys/0MlIDyHs3AeoApgOhZs1FC
pIuNbK3NTEFwTk2PTNCzVwUmWwb0dxIsNhlHtgCH45CyP4OyqHdHMkoqrsUa4ynvgWP1gDNjNZoc
7pPEsWfA7TNI0WOvf1mmpwymtOkOrFj2/0GzKWVxQdWmMjz8GQ9hT1E132lS9dyHU027cBVnQaOq
UxL2sToR3PhO+eYpq0u8Hm3xKCsUcuwx52mLWcoUM3SL6fN6aT+cwcsLhuG3cKkQxbU0qm2505ZO
vkc7on70kZQW5ErrsNZ7F3g5ODPwLaN1/aCYrb3+JnlzFX7sNZVqVHlCncExpvZyVsfBZH8mWApG
OWhBGjmyTwvd7RkYDD1gJcNF9N2VuItO2bZwG7/sYfZjH6rA8wGBWbBt1w0p/0nbVV7Ub9hYlJBk
NkBMsceevJquCuVjFPJAnKRPCWSiZjdiOtzw6wHXT1TZYn4iANo97GcP4PYedLYjp7Cyz9XFie5N
EH3tcilQrTE3A7MttFPH+Zw4DinX3t57dMfFVWAVodu+FmihKYrqZH95ihiE1hJe84fd2rd7N3KB
Li196q+fikzUCuaV8wyETa3gpVtFaYtxHElMwfgmtev2qUzfqZQbVoS95NiWpNIMHbMzLDeLFuGq
9hYCBVFIwl06k+G4FP+lcTaEZ9B8KFtzjazw5dMBh/q6b+4Z9xwrIwHBUzTG1I1H70NvT67tCsuz
HtJQJy1etOlErzuvXAUHuyxADfpJHxaqlpdIc01NrwbmEPwLJbscpSD2Pvvf2aKf1i/0yfzBVSxB
CvH3C1n7j5ilf8zhQ39cAMZczuV+aKKZxBNGi1ml+uJikZMw2gCWtrKaGaaHQE4byd6qdYi2410d
L2Ur6wxQv3Dv4bGVgh5M7+ys9Q0LunRlvseToLhj+spig9fowYiQukKuOHpvaMmrQ08ayj+saT2X
WNiYlMWVVyXA/1zR75FLVSH/4XPrmp4wQUoDYtVl2/XW9XYq0LhhRppwisg+EzMV09YRqmfFdx00
tuKskPcXFMVCC1Mt/S/Re4wOGmHWprNisX5oRbASbctmnp6Fq97d/gAj9SR/ZjdL2QTkrKSuqiEY
pno2uSXG+VsY9jednKTqOurc4whg4kdzWiTsdrawoSegA33nMoU/1bq68305mCDlX1G6MwFl2q+i
FBPMCK2+k9GA4uC7J1R/+Lih6lotHT7AmsEeq3ZWyg2Bye09yKf/SBnFXk/8C/Srfni5B6Aevz9o
hopzo1obyyC/wM3kvzj44Lxq2x0ZAFc/m0Jj2kNV9SmLg3llTyObfv/dS+vQq5Xiyj3uAFLn3t1i
xo9txgo7Svrv0dLNSWLkuGm3VEUUq6jiPU0uhNdlPqKPTnjKbsh8TGMCz7raBbLTfFxGno5fNQBO
dyRHg1zwyp0adC594oJErEfhYCX4NRTXSHvLbjQplgH4BdDpuJmatX945zkdkMOx7nfu64vY2kvm
Av1DUgL4txEHWDznkbfUXdj2QIe3JsOtmpdrEDu9NL54+QbH2P2rzoqH9W0MQ1dNm8rmHZ9zMr4L
tpRpOnRfirooefS6fkyiKgBJzyy0oYcNWrrIt3kmKU4cJUjJlhIgRDz88Nu7HnbugAnHVi2uJp3O
sA4xKVN5sEJs143F2umdY5WLLIHjj4teCs8rJg2iUrd/X2mxMB0RY59efJ12MfopBGoX3fTPf+vm
BasHa1r+aOOLuSjaVQeApU+9aptd2fyw+L61XFJcGcbH83FMiGxX3oAB0j+uUVwxnEId8uzVTBRU
EN2r8u5cliO4JnUeHpBmIkWMtXkoKbOJPKtJ59Cijky5ANITGxQdIiigkjIdmxPpKRkBKshm8THs
Dass+BWRmm2ZnAsg2A1hvTqRxKexJh0Nqzp3vJHpubuv+39P6HsB14gSoOXGxdHkqp5Az+dolczp
MCEzCekT7mt7shTQWiUg7tsj1KCKafplrZPY+lvUz3TrkudtJ7WuBZ3w/dPGkh7j5Pl20Sx8F6tY
ujdDVC5U8XeNRlgrPl3QkGgLIVI/VikEph13LcjsivmUj+RENf7BsFs5Plkt6pv6/TpTm/1DSXN9
CLs5srQ2sT08Y8ajzJOR81p0AbUI9wKeErPqldmfKC22ajslFirZylerVuZLxUzqx2WUtXNyykXg
two27O8CJX4LcPeaxrTE4uojjtZw/tKUBcLdJ5WajHZAmZdzVeK8nak5gbXhd6fJFDOATcOYWF0o
jm+L/flxyTxMB9/dxWQa6ZNHEtobcVzM0gwY5byT9b3RN6OUdE8j2NaGeCA4HAORPxzhF0lN40wd
2rfPuH/4ykM5gtZFlWbk04d1CjRvekqvoGsM8Yh1BdOwA6ekTvXxTYxOoaH38jSWFDxeOfck5uua
4XGt9wYvTTv3PA8pb0aBFWCNB3w4mhVpMHPPIOxLBXwkCA0sROSUxC8xx4T4qOaW157w0VL6SF/8
4mhMHU9RYMT11A3EWS32rvVAS+kSr+lljUvmXHqI4+8sRgbTo6gfXNwL4ehchR27f1J9p3IlrLin
pUeJPb4rR+mJziPTLvoMA7TZ7Hkmgj8p1dA0Ag/y3k7rH8AvJwbMvtdHbt6Lfc1k5wkwlRQLQ5Vd
xTlKCYYb4qbKjNGaLYtxP+SROzx5advxbWDksyJ8whKy0GB8wQdhzOnoWVKGg+zUXm5hZ/exC2sI
/b6mvybjjMAR7uImYxGyzRxxiu5ggzkTzStG5CrJCUKT09HlglAcRGUecc1S7Lfzp46q7SqMoOfd
Acow65KCLJ1LkMSNANiu46ZhdDYT9maoNTPmHZOGM/isclWqebgkcN60ipBa6n7qfGZSgQAHlXc0
337LaXZga2+Buy+GmcvleRT+sy9QRw6vzzorQu1A7oTcR/Cp1hr3oYiiDqVQqqUTLrKhyxtGAN1S
jmSoewW0kLTB3FbE/wkv3B0C7uhEl4TBqwnKFAzz4x5/7D1sgel8tQf+0RsDoyb8bEg6lj5ZLWzh
P7o0YiiSEQeDier8/tMBM+7ZL0UY1BNjpdAiVrr3te+yaxnvi8dc+gkQ0GoZbq6xApsc0vFYbljZ
hUL6spufN2Pygy9tw27j5Jf/DQLcQHtp8aJv71YRiucRerxdnr8ZO7Cuim5Qg4P34Zm5tN/ntgxz
IxiDD8+kwBDD3BLrD3C9UQrVsAXT7cq0FjQ1h3277x6Z6o5WZMXhgg4mNbyolb7BfFtifCpBhbLn
KQUslX860PXB9wkjffOXdbR4q4hq+QjQUN1WM0MSe3jHOlvAa9au3XfCH99GQT+japqHO4q35G1p
D/xZu3rasQAdlkoH/LDVROAP61b0COSUcYnXQLqILoxe6zNHE3HzJdklCwTkJ6394oOh1ZbC6x+U
Fr1627uOQVNZzBp/l/Xl0flKA/wfuR9jueDCstiSiSg4aymgBHZQunx2qkH4rw+ptkWgQZzcTtDO
1aEZLIKmi63NZfWR55gzPaaQOqLUvGaPlp5rbagHz5j3HDP04sx+QW1Ln9MD8p2WnZhI0fWizV7x
gvtML67hkmpJZJkf2JN33/7xgySX4IhvrdHmB/Tet1mwAtNpCA/kN+eFWS1jlv4oH0w3IEdkUsBP
rUYAEcUibKf6z6bt4o4BIbj7Vk/GC2lfKdGwdhE6ZAFipCwAqaAGUYCJI80qmBHBu1XSn9zEvadr
K0E146cX4LnM4GmNp9wSDS9MxhwipG9mWlrlTWP9UNgsb4c9XflkvjuaIHZqWou09yN3GZWLJ9gw
Q36+cae/+VCi8BakZGqWxI4Lz+cYMzZKpMPnoYSiMSLvKyBXW+bH2is3duRMXhzMWW84eceEEbEn
vY2vtYq2d5G+udFMlq5JadwkDPIPhTcfx447v+oAbxxLMlXlm1QPhXth3/P6p53deyiCxbZrNhT0
Nje6Qo3bYxek71ZVADZ8wQrl18cQ2itEJxcoU1MiYHYm2jMGC45fUZeEeP5jMYVTkzHTi8HteH/E
ghUj0LPLAuPOJp1zVlTdyLFeZj4M3X5g7IVeXRpM+MFB7JPLuRHLlVhwxGsJrx0ZUmCnKF1dNDGL
Og1XfMdi5mqOgBh8k71njZAMVpJ0Hdij94bhb4KZxKkXjecjR4+ja3tPTuM5Lh3LqaAu9dNQlg+z
32TOCS7+oDytg+FJSbRAN86ymFZAAfmE72lxbOWvRU9Qkmm74KV01OtRS0jFyXUP+4xwXs7jmsWe
XyxjNq2NouD2vscVeL6jEUSfEtor09UDe+ydgZ2M6pyciMcITzPsDir3VRMxZqc4DLYxjRnEA61/
4+2NfF0WPX7nDbdJCsXbHxWD9HxKxRoCwkvTbYbYZRTM4TlhvxnMWJhM0NeOfMp/GbYHEeT5CqHV
Xze5fYZHs0Ls7XNeX7ChuNumKK4+GseyOIxtDW1gx5LDV/np+sc2D6JKzHPp2E0/cba9BL1K8MGV
/lZz2ijqtkHIKa39DtqCSfGKATs0yP8NZ4aB1CsBSO93wSAOMq/f4pzprK79GCkSuy+bZrggI0iF
7lyY38oYbtIkuvMQtMEYQ+Ff9kOPaGETabKYMx8dEnEMZoq649SZNLH0SKnLaF3iDzpN/mNZkhc9
SKU9F0uhx8qUSyko/Vpioe/W81aHooJBfTWecQvhicPZ7QNNHCaLgNr7z72aThk9KpeOLcf9Tu0r
1t81Ig5hhR/FfGOVde2B9zHJIzkNYiA70AXFFMxPg3xjD0KRFO1KEH6stP/6pnQkVBcq53J8Bb/B
HvYwIf170vvH3mPqdv6Tq47Ns49Mtpf+YOzeXlmKZSUSBwLQkmSfsLA/5DDln3oKdeyqhu1RoW3e
/K8Dz3XJnhpST75tJ5F7flZjG7EXfXl0scc9U63yJLRZGavlARgCrx6PL+lmxZaN7pj6DDe2Qxi3
ZunKc5Hkg17hiPfmjr6CIbkIIwbEsVLLT6oVo8RDOoL4A+Ck9eFHUcC/NkM9mWluXMVZGWvdKrcf
5titsRVjSOJpIDJqMp2dZc+/mxq87UF2QeXFS4g3kihBKOVejXt3cvZisUMFzGHu8OiugVNPGkYF
k34Ns9PtZIwj/iuYqhQ+OgdZhN3XTrJG/qPLXmog0lZE5nevxJDbf/XbvJSHE1iNkoWmsYEcr/AT
6VZI+nvIGQIIusiQy0ot0V/2h/WH8EwrLy6eZnZha4+KqYueK2KlsTELCvMeG9dx/5jH0W41FEfW
m6CbxdrjNpHVsPyyJ2MYN8/tmf4l88brM7f/7V1Z7XqOqsH2Av+1lOg+INcfGkTVenilkH0pATVz
25zsyBYQopV91+JSP/eoVEQ7QbTGCf5PLzsyPmfE7yMMiuJc27NgMsVQuziUjOP8AEM+oOEPGBlC
N6xZhWVKhb9QzxnXucVYb1OAA8z+0TAh8PbQ0qjW7hr4ZXYh69Pr0zdXZ5JluR2cBBxqy0MHLzN7
85/Heju9gDPNzgw/9qQ6lHDKWTLzywDaNlE5XuKzdNyKl2MpgBVet3WDgptkUAhT09XbvrMUqtb+
PBLYIa3CQfAG/D5ueV2bIrDW2c5c1XCMjxJQBYAYqxRihiego1Pk7YakoVixyBP9mOiQF4DZjBNE
auy0Bjw2SRlJU9cJj7e89jA8jODi0LNys/btLUNsMlkKh3ySqBZMte75vNMDcZ0SHsv8R6pdPSFG
I428mFFhQTS8R4rY/gnSeTizaRbrOqbyMRqHNuCOz/3BudyJbVl6TS97ApwEXY56bI57N8ghF5TM
U+Qcg3NR6nLl+lOQSNfJQTRCztY55rOOBTkSxEdpJo4HKGTWE6/5nq2wHATFejyLoy2KdVziE06b
4UGxAeogbS+dfAlc5Jjd5V9Pw1IRw+H3yMMI5SooNWIn403qQFzRI8RbDOmkEbTgFFq/V+we13p4
14CfIUWmrO7ImU6AluEc3lWpt+t9gqJGBqeONDDpxR7M8KfMeGk3oEcLolt4POBwnRoP60jrDnn+
CrXsU7TP5qWtP/rz9wvuSSUWjXD8KBM4n60ePqqK3nNCcJs+cWOOxl3WtzblESQGTDKTqm090FZJ
IB6kAnXqGPUnbjPsMuqzbmjBfzFfZlM7M+L2fSCWPGcBpz29jIbZNopDHrxWB3n5l3XuyoKsr1bj
go6/RgyOMqjyVhowzHcFjX+WPwRHVJzYA1L7jG4uG5OVTaHWOii9jpNHtIqcpoZFh2vVFyMj8/pe
yh+iqYUCsvJ27by28DVJcCJ7V2XbNAN5Pq9aXPvrBRYCcneK8TjWHBeUalQxsRUADQu+6itDP0w3
VNLfjlc3EpKUoA02ssZax49v4MtMutK+4Ont+XVGIv8rmcTwrMqH2Zin0b8RwGl3KERqfTVBxiW1
JviANuHYbASEwyrbtRHaaEgPvDbl8LOOq+RbgQGxxunqRLVdoIy9wZGwXO2u3dNfbmgmtZ3w0JuC
2E9E2WO0VBjQaL0f2r7U8yz6r2WmVDKjKhXMWsfmirNylRR/p9elB4D38mNS9YlAAMp6vrR20rHJ
d48Tca9n1wPj5pJNO6918166r88mAjXEOmEhwWmAAWnkU5PiXd0F69ABw59XlWnTyCEt7VtrtuaD
RGjZRQf2PHEo8fCx469hdrddzY1Ewq5H0pCFeUXZVLF7EIhisJhVlZ+QHDPomqIE3TGHV4jpnZyu
JnGMDaJDGGrcBBVYAKn0wvybt2Kn/H+Seoy/gbmCHFAzT3ru4AhiiLhA4iC5pHz96WoB2VGvpt0P
BsDiVpXlikxMT9mHtJVhAPU3buTzb7MR2jj+trBst46RwfDreoTmXCKp/LfZqrD9+hyTo5KEMNR+
OlQ8mm/ZiKlX39pVe6+Km+2XigZUdiP/NnLMCSj87eJIAozR5Y0VmRVJ6iuwZHgOeVYXZTtGAq6L
hhcT6Qnq+bSsUaCaPwOv+QcScq/nLGaqTpV1nE5jLmEmpcEn8DQiWHC+o/WQ/TE6orf181uOreTK
PucLEpe66dFaZ3Hq2Q9qs0AUOVn4bsaMIlHIvCaF5zFTFpnVG5PyruYJLTUH18DQw+D6+a5iTK7K
kvjdfDC3NBP8A5/blna+YFnjTmzypYG/w4tKmbbrK0iVK5L4xh45JUhjSyNIUeKjTOZIk/pkmSS/
AbiqQuJFMx+anJDdRns+43JyZAfW6rPLuft86WRdhQdx9SMFDe9c+FUPFjph2sW7ldraR6eejVNz
dZj7Aw9JZwkQs352aDyCbvQVwIUpQa8q1f6Bad3fvEog4r6EY8dRdmTZwJKIMhP0N4G3PN+z3iP3
9Z2+ym7BFMPb27MXyWrpE5W1iy+LdhOPD4NeP8JsmhQSs98nIJj5isSScAvZpoSbTvZDa34hHk0V
Ko1CnoDjCYfeeKpmDqMjDbej7ndA8B6nzTSnU7sbkSXlKWxRj0RkEmtZgmQvz4PzGzFLVwO4WmQm
d0bxwY5zXJskd8K4Ea2bUYl2geLZjAx2F/riZLml8a0SOUqmdAd6TNpelp2dpwuSTgJzIhUAzfbW
utEivuoEEV1YHfCTFKt+KJ5pXtSdpFFaPj7KJtEZq6sxVCautAh1RjvtsFgeOUy16A5QocAsra5H
soML4LBNwg4lmgQkEZyE/x69xNp0wa9mMEYbtxcQmILmT/2k3EfE1/2GOkpsj/VN+28P6ll8bHsn
y6WTuImma9lSQkznBLrX8TKa8lXbzMt7kcckFXiHbqnauLo17Wacl+5JsRDXjcOF5W0UYBGnIvIs
zUd7TtPF0f07eDjmUnrmnGUNoGzwzFJBPaDk1zS1dYtg/Foy5lgSIcpTBLu9q8C2scw31QiNQich
bRu0w+qYyDv0DGKfAP3sxMRkbIqn7qfCmQ9l4j5+3n5lz46KQxNVcrbSJgBjLYVd0V9uTiQpf77v
4y9MwqmtuKoQu5Q0vUZv+tJ4r5FwImcftMAefjpLAO9RRjkYa2qSnsQgwv3pMIvazi8GH8D0P74c
GYd6VS56dfuGpKPELc7uCn/1RhvKDdWXWnfJZAvLkCy6rQNtCKHtjqESx369mDz98ou/PV1u904O
JV48TOqrZwVnXu7mLrQm2x4UiRLU5qQ7/Gwr1DbVgQBvD0MuXFNhCUuT4yB+zTVZdRHO18yIpEVM
yolH3+vOPvAAXvJMpgzne17Vo8ydV/5TiYr9Jb/gXDNpOQLTgYRyjh0vHzBSiAQi+D4t72fPFCeI
aug94qZgQIUgNqKfvdfv4RHrBZT5Bm2EE8MkBiwS+P++t96xHBl1dsRwLMjLfeAwowSNba5v++Jv
M0GO91HgAuCS1whBLUYTXkxw/k8y8De1j7gBPiyyvLC6fZ94nqBE1J+jGWTGAoMkG1+cp31KBk/U
LbtDfC9675rQDBOfnc0G0X0X7Gia+HzIyy1tldqlHlgb/7VQH4Mx55JXE5hmJ1k7gLs5FN14jXRw
h2zmhaAz5vnTAvJEVakvJngKO9StxV2Jan3ZQ2uNWesJN5v/uGbvInU03Gt0Nrba5nsLJB5uo604
VP6VlANqa3BWXpveBtetecsOJBRAQWvm6hkkL/FCxwsVWuNsztESmKmRO90u4PFRyp1SFe1Ax11z
LfOr2gRVSXqADkImetdYzMCNo5MnM89uycYlvWjbGnVSRINgK5WdPwFFvqJh8tBuhMuKpi8ic+XG
sWLPDWzYpwCI/lGt1R4mTzCxkWaVCc6kY2G/1StrWqXqPIVkgmvgOayPDg5QMlgrtbpCOa9YDdbt
I5o0vVGLcz/qyeWm2WxF+29KImcH+Ax90gv+uBaibmiwH21B1hu3kJ0mgvTJu1LHa0Lk8i3A7Bvm
uS96DmXlZwD2gClKWl1OHc+aOYctVPpmKvcYVHoywoEO3Gn7zSQss+UrVJNFSlJ4Gu6RZwFtAQO+
wGtOHSlmMFBats/PS2L8pZg2w5XTLnJbMaSinsyV6WfUTGaw1Lo73z66Rnam60H6Dbs5Vgrdg6yE
srGuO+WMDkMKg7lKqryROd0LJl6+3JgB+RSxq1Av2eEVz975XG4gRCJJ9rpTvbj+9MnMRKGZsYrj
6KEcuyKnyYpjqIA44O5xmIoRRcUGaTKofrx9fmVe+hoHLVaUsnbTXlKbbfsXgaRz/hYawgjb7Axs
e1tyNGRtiQsYGd7oSIWXAK64rWKBuWNHHtIQJut8GXaGBzS0qxtZkR6R7OBT0G63hUqiH1YYXLWY
r0wIDTp4FH7OjiM8JRlvHwUlcBMA78htYlH4t83WFvN1Qle+aEq+0jMI3Q7YXC8IvjioLzcNn7UT
5UsUn/saG8zHRC46fzRuLLWkMIvt0bn0iH0UbeSLgXHPCQHS6aPtDC82Yyuq2JImzmQaRsjOQ/rp
TjQURt9WjQUpLeFtuIPxbLYXu8PwFIg9wEbmRvip9AmYEHU6yo3P5g1ZgaoLnBFwMHq2uTID44vi
gC5K4B4hNEG6px8sb9juvHegMkGKSsdBKl8yOk737A1hJuZgyQHO0svKZ3pg+Wce8BKQArqMX6da
D6c1q6sarHJJIA8Bfi/q+yNaohepfOGEOFtxJH+ClDiLW+NIy+jRwsJhP7mCQd1KEmEAnKE+SBwb
jSR6F8LLmNH+0j6T2e8RTRDVPD3P0j7EwhQEM6E9URpTdkWqd0snjKVNms7TamPERDyftAcXmMxc
s6NEcXnVWhKPpU/nbqKaMDhoxu5rLNNXzxlGMtUmsCq3T6atPS/cuMfMjBwNc4bU1jSQbXKQa4if
idzK3DIw230PrxlehE66TDOi7rROH8wYbZ2hjhLtZI0JiHVL8toSvuaqbLmrT9mg5I++MZZGQ9BO
EI6u8/aq7i/J4Eq/jFgeZLpgDlNNnuOBel9Xuf/nM0J1kNywWV+GeuRQXupy2jVjs8QV62YfWoXn
6VA9VDWqKMMRYRqvN5C58T3J64I39zb7ibC0AMPdYflCZO7DKkpss1ZJAtvy6jkGk6dGlcoMlCAX
nY+LE7J5BVMw/kDCFQfea+9uLZTNlaS2Ee3lm4z2uPb5FaCoBii2Hiwglyt0VL9at65dAMlGaUwi
pYYC9cWa/55NY255eHODxHSItBMOzJjwmsuOOAb9sYZgxBBLHui4/KM4SBjpJmRWYb5bIfR2RKdG
OcdFi/VwtwA6ZR0nwgCUEBRq2TPhqfVTfsoGKaykz+es0CrKVtQ4PVNBn/AeA4BWqXmAQ3Qkk0u4
3gnHm1oeCBBk5LcRs9KTnqwlmNVjS92r8qJjIlq6yTc0CoJf6rmE+16caGSMH3LduBonczWgr5aL
qsHAvJNtWKHZVEu4xThdBtHNj20BZopF5eW1iPsYv2x7EDAovBVEKdVqWvVVIUdBjRNegcKdMZhs
uRdtMtBeba921tajc5RPkSUKGQ8WMQv6nx6VKu3lkfBedhysIpam72L5NAwqkNoapZFXq9Nd23wL
GrG66Ay8mz0qVcspV6CM18AlmwApOeFRZe5v/xAZ3IJdfeTnqfJ0bsYj20+KqTO1KoFOGstpDBri
EeJfZLXHQPl7TNvl780iopiHcdvih6WaHRHhlAFlmjWC/RCWIqKQVp4r0HRgoWbKZa9KZjp0nRTu
netvbJjLOxtPkMjyTt/C3pKj+AeRzmYg76zuQdc5oLoY+yorCy8sNjaTe3osd5OC90jelX+1DaZM
Tnf2OgNLqkwqpp926JvgTCl2I7/VChfrn6DH91rXQeKFujmwGAadvdhWZAcNTWMtyz+3ld4DdIEJ
bKjZTPd+fK1sVHiKNLsJp5bh3EKFx4VpJGKoV0gX9YNlrig0MegvY3wbwwkDEfWARDlvHczqEiFo
T/KKvkHmtz2o34BeAvGs53+OChzQpkR8xogKuHvQ4AOdSylcpwcuUzlR+JVUUeJq4y5PIsHiF6WJ
OSi2iMSucR7iabFS4aQKxT2B2IPsIdxZE3aokVMZ4M9jXbf9cn+5sret25Bu2wSJimXXlBK99k96
bIPtNz9J44gly8DuPyNxiuotNkx4sKVtJ4MWeelV94IcJbG751ZtkTsENiZTdE7BMU5ZW6TolPaa
z/0M1fYLNUOu8Gm3ARMRHZoBVT4G4WNr7ddNIufDP/ygGbCarJ5eYT29lH3/mxXjuKucCXc6/kC3
ZXFgh/bawLEtV1fa5P1iCPT5qUxr0jtnxQs4IJzA0MTnhUdKxyQQJfo58wp01GAvICmKP650XaqP
ZmjKnEMjLkqPoPwXTbdybO6iVtbHBPVBTBPvRGth5nnK34c6KC4y2E13y/vAsdRGl19SPAqVrWO4
CiG1Yog8k28sRpcroivAwpC7e5vyPVV1Q/BuSAuftZnOO4Q/YglecOOJXzTd/LhEVQS0UXWo/OTH
mWDXVbOxAmvOE32HEDmdTLgvbmoeAeISLAwwePeXKrkHnn0X3Uqapm0UgmyaVkV7Az/0UoxveYE8
Siik/1rJTz90ocZC9V0mNFO/gtyqxfgonjljqbgJvP0PybBy5cc7tA6O6QjvpsfI0MZHxsWHYjg6
sz7Tc8TsYYfxmmZ5P7UZK3YPJqhX0ppH5VMqO+24HRVlMd3+PtZHohDgHvSrK4AmjTBptOAt8hZi
lTYhHMUD5Bm9x9t0hFbwHyWbPnfnvUWtc93oQ5CZ1B9fZihS5zCliWqQbordtngzTeUxdTJCSaCW
5vJJ+VoRKCT97jWsAA47YKt0wM5dC1S8kEgzZpBndCttaa19b+bG6vhCXq9a+G4GTImtmKBehnA9
/AIuY2VlEpFOXPzToaz1nnvd97YfMzdXzc/EqNv4/Qoiw+3WzGaB9q4RKiKh023t52RcpgAExcr8
tq4BqZGLodwj8mMbBynAVBcTEQ5SBeu6AF+y9Vg8xzDCpgGBwD3UlFPki3n9B0ss6WzA/42jULME
eoFjLje3qB57fidIayxRjlDBj/A5oG0aIn4kM5Sua5cs80bBlzJTdwEo/KNw4R7k/4pyMxczbUyC
Ky+KqBvkAatirK2pNqRjjYStxYWERIs4sr5nXEg8DhctYyt5c/FyHcTf99iX7XzPgEIrMIDAxCvL
yXIuwI7lDAGwnL2xP5yiCVjBs6CqHKW9HLx8bq8ycm24aAYdar5/3hxhCrEpl/kVHtUVPMGmUx10
s/xPYps7qeK9wrJO2FAfDluIFwTiMYHa5wnVR8ioK66BcbudyljA6R0xCRzg1cS3DvwqCNdflQqE
NeH74BM+BnWozmNPD3HCg+Ha0Dzw4ZADN9JUEr3hOoO1qdUf40l3yBaUsIFmAJQ/PfGgZVpbnu1O
aeOIYkX8CpdQy7EBmdkSlyqFwJxtRs34Wk6ttj5w0vkuybsuNSKoYS7dT7p1JGdTu8id+36sZBB+
ZeCly8E2b2aDNW3/OSB8DTCqAl6rI4fXknS+/vC5oWyJyuDwxYV++D2BZdEXntHizlVLnjHYAt6+
bEc+YzKCweLX+/wydZtxrT02axqoAQBNS5tPmnA5oq5xTAm4tLBKtOMrBsgiO604ZIBJ3Pdkd7nq
gQZ3B9l+F6BKU8rF2Dp2dDnubXXpct+kYeNFnrDQZjzrN4WBzbn+p8KEXL7bK0UE45lLEgHYV9VU
/oR2pKiQYppijX0lPf0UCbM9/WCk/rECbWJedoIljgjeb6l2rL5FiNq1F8GpIeZBNkKVX/HeSv+S
i2+7ggn+gTTTWydDs6OtPbBGIwN2d21ZUpp+mXmN7d83QahkR2bhXAEb/y6OfgXRLtgJEX0bfTQJ
Tq2UzgxK7MqknRvg/v4tQNXLACPMljnv3rFBuoNgr5nu3ccNM1Xqty3JdOanw7SWV+EpNewxN9Wf
W/71q6ssMWeO5+zjuCSgroZJsYoTv++YhnYOX9kXDbB8YLRDrHRsfO7mQOH5Du7hlHEwEhtvgyWM
Q+2n6YGMDjgh7Zap8V2bdGhabIWGAsG+3bJzG7imLUl2fnfLONqdKSxUXiaOfvuLYaJY9bmolU6f
JCpMMg1PX4iPW8q0sxxEWP2Q8IqJr4YR22hltCL58TpAapMfdAPhsBcO4Y8SDhSMER3c10J7aNFl
pcW1aS2SUAEupYDtteacTgwxYR4hxmvOi7XbCUwyWJJpYNDly/zNhS0kswoWEF649P/IKav4+5Hl
mPVBGTKNnrR3DqU2enktIfDubWrKs0fqq0N12zAZiS4fCotBJfK28tTpjvEO+BobTD/lZdzUdyeX
WdF+TsjOeOgtCtTtn9Oj5ek54Vtt1TQPXxiQh2Nqm0fB0d6P3Sb4ktj6plMovoziNvZy4mE9hOrg
C+NlBHf2pL+yJxuz2/sd+BcgZ8y8vHfoebM0UHyc2CKhptZlRiuvhmymjabKN2pOJusj6RTQ7qxX
so1B8+1JxSsyCZ05NXTPScUDPH2bBItsW4K6kSdiVS/spORKfrgqmwXAjld52FopGk54WvNUlO+M
Hk5plfl8LwYZ1anIxqkULwZ7ZXG+pkaxWcg4UlKbD1PLZVnn3CHvEuxjfBjvmVpsHRimKuAxSjde
8FpK7RERwEeH+KEpL3Y062NxdCPKjLjoFusZX9t9jKgBHiqE2oUbA+oux/aIBBvPd0+3HedmVqte
uuXDmIsOa+zGp4KU1mFd7kCyfb6FQVsi2rwphmNxICyeW9p2h5fxn3aniYROQMUINKALocUWjMwu
SnblurspqzEoC8HxICXK+1Sz4hEG8BQ5AP7XW6tCQCWU/tdqL65p6POJxHp/Zqa1iamlvX7aTRUz
bn+iCDxMCUTd7/OTI3uXm5/XZsjeWXoTGHbeU9JSYCIZyqfv6J/kIOnXrLrsC1Zh0a+UUNYLadcE
WhmipGy1I+maSuSu42Df4RUqNgDvc1uqzOMprCI+S+5WU0wKvld4VmwkSIoZPlU/CQIGY7kjKfJz
uMBbhkYr2aWJDMahsAr5wwMH5V/QZ8RyndLposQ7BPeCrHGjP5t5tgYCdohbeRgmt2zx4FO/lGDK
G48OPPOtw3KHIy5p0ISFVBtmMakUS/oTu0bqF+Ouj8xihh4VJfktM63LBx6poJ3YCiNCfSi/3Mwj
NIrbESo0kxa+kGN66cHzx+JXLjwcE0P03VOZiP7DwODEYC9j8lSUUHOfAniio871GnK/p5JyU026
E81pCmLQ66PEo7MTinNPE5uZwKw8st63yHjj/YkpbGaey+vUPOCosf4Oc5Z88EYRDC0rFxJNuw2V
WNLpirQy2FzNAFVCHpMrXweupS1cpoxE+pD7aFzbOKbbs/XEgjF50I4w7L6tGwprpk/44vtg8ydo
l5p/wcm96VV02cEhHEtZ60Ica2xjaysKXJmSG2JkorIAfN0s5EQ1bsXmcfHq9wnWlcuwo0OBO7oz
AFuNvekrEkFFQC592rz8vnq4Og4mdr0SR54YTKHFJcqJYI1cqD3cYDD7IaFrf14veuG+NZdZI8um
LyMDdRmCN4IBK4Ci3+xOApGG0F1eSJloPR26q/Yx+1Q/cOUAv102Fr1mJ6Zxq+mXT2XyDUtfNO0D
S+z/l4s6Dt8L8A44HkDWaD37RVR5lnItpH1+YrQSKJnvJ5l/UMe/AalexnbQvoIKDB5QQ8p8MEGf
wJWGQmTjkNcvhLf8IcMPVEfkA08iEzXTWmDWTu47TFu9xlUjSf7gJXq6XsAC1kw1+gRRHWr/PzGj
3/1ls0mj/dg3ihWdPLFJZWwQwJ/RsdGsx2POL+PnSn7idlaZCzu044KUSQ24WNTDYUwu5Bt9xm7f
7/pG8XLnXdzvqZdNt1UHCaHY9vI4jS+3YHqjkkEBXTEqx0aCLA1NFjuDAriyWZXXZ4GtCARESirZ
1VbRYEH5pOmf4XUyNKShf4IEU3Af+W45xnob02aLGZHtNB2ozjRQOOHNJsoaJJTqoxoOORxMUS4T
MBzgHfMZccq7KyjFluEjCBSTKx3WX1k9gGfCg0c64mAnq6g6dHcse/jugJrao7XFZowWvs3KiE/P
Ztnt0yufJED+dh5pznzrZWzBVSvzABSD4nmo6Imaw5OyNZJJ2v0pDK3BVbgHjq9jTnAGmnvOi0D3
EUmSRiRYnS0JF88vpZZ8zaF0IMPnIywZ2QYUaD2JNRNVwB5mh5oqT7l2Nc2HKaDbY1fHWT2KP8nf
uFUvU0qUCU4WI17SEvdSkn/T0bbq505J50fNEW9UnvLzyzgq8ZIZ6/Vpu3PQeuvWLoPpcmRbsJW3
BO6gKyI9C+tKNNwKfZ8DE7C0VLfSpmp+DCi+pJ4deWpU3dfmmLI//eZrM8f+0UxK1eu/F0xRTvwg
wpiKUPkV7KOSuewTBsYnQqTwRHfyq9XfnXW0KquaWoiXFLDTg3S7XXQXN6WuRDEV6MSzJIG0/FlF
+o7lXL3o/vDgal3KsjTvE9r8myqUVsI06UbS13oO6f3oH/V7m0Zw1qO3GmKxpnSZBNj/K1JGBYvY
c7oy/ZQwSoCtUotJHwl10i1S5IS7aChmdgqCRsq2fEnn3CZNLH8GNIMvDAiBeeGhd4RRm4pFFU9u
7UbzS0AZR1uSHgxld1Ixl0M+Wbwl2xKlYPwaJGRd6BBlsb9ZGPUIClRziwxRs7hP/J7Cuc80ma5W
MKaPur+yfBmGWJxochYRLPzN1FfCLWBBz4pq5DL3cSnSlhH3SHJzmAVZs44GtFGiId8Hx0DObiWt
L28hoovyLG24k5VG2IO6J9C9e8QIheunGqHIFuHrqf4X9y/7T40glR8b1Pwjt/3lo61csC4uFzG2
HQ2xxfTfPZbdLc+8kuE3W7I87Ih8lvMub1GGLaRCO79xtlgJFQT6Xcd9n/DpRRUqxReGsW+iCc75
u+9Bq+wloAWSQz1liudEyH6f/sAhEobDV4fLMpSIoFHHOS3ZvaCTJ2a41znomSMQXDthNtDp0FiR
psBptxBwljxg4AY7qObgXJhl8w04Ts4zCxvZc4Kdhvt/jQzVMwPQ6qcKQ6XI3f15Ul6XjIVhg/qu
GvOLbOZZuTnN9JGTXxZPYIdC94z3UySKESIgHyTQfvO+b8kaaPWWisnBglCgBLQy3GndMJYFfJ7H
1TA8TNk/HOiGrkcO6gZLCLdTZlQfD6P1xj6/MPz1FY5HaoTHxK2aAxE2CRXcEgFUdL+S94YZAJSN
EWozlBo8rmuY38lWsfEqX53UpSruGq+ieP21JE/Qg/HCWXBMf7A4FVkEJ6Xvf7RnyWLNlyP9zSID
RwoEA7I6n0tCcnFnzMgTBbn06h3TkVcP15DO44fGbD8nhz1N/MqLNur7Acp+yJ3eNoLtPyc7Ujdc
OqwO4IvxGtJ1Lp+5aHeZFURLVOSr64RJnKmNSxYi4Gl+E3uQ2NhqowmfP2kDZWdFTNvlSXsz83iZ
+979gGW7n7l1S7M93iMuJR0kE5KDXgLqAEJ49BwB0ytrrj4V5kGHIXVURyJvpZoU5nDaoK/gn1CF
dGzZbLPWXJZtMy/wFOUjQVzTr/F2B7ikio7SQ0M2iJ5tgQEXovWQ7K/HhBWPpMVZKZBoNXFnp24w
JM/4HpSDuvdxIvvIwhZIPddc4tivwMC/81j4pZf1dvxYbfdf1sDS6EUXUAQ8hJovPHV387z2Gqrb
K35snhx/Ce6tOt5dBYH5U8/ETAKSUXRQ4g8GMGnuQJWu7YQlrLQo0gMimtyEENetohXhVtaAj3Of
oAgZpC+C5smkKum9EPuQWqgBJDeGNp+fnIJMk0Qpa0MeCFw0/t2/UlpJ0MUFAsghbdOSFnnXh/15
CXajwQIT20D24cWh/OMQcUU1u+hp/dGsvXrqVWYMN2NvmnWXTVebOSOXMaPAiKxhf8UTuKdAAYdr
V6kSx7qULSGvnUqBtYQGVUMW8FckNgrd5lgDU/59ZUfV+084alIX6Y8yJtAdh5QlYaCc7GYTCehF
ETumUgARdKx4JLcKTX2p8WqyaEmYM4pfJd2aioJ/c1+T5pMq8QKjLivvnTUZqtSo/dhxyDFZPJM/
6Dxxjhp+XA84C2ZeUAE9nyGZuFn0CmWYEfNU+YdCXDeUsia+1r/2+ga1HDDNNwGdvde1ZgS5QfGr
k2wEpeW+vjAw8zbSsnY0FYDHKC5OfgTktva9+eD8Y1VSwtvIvHRZWEFhn7IIFeOz0gfaIMRU1Rdk
6yD46NWxs2nN6jNkolPzzNngiYe5TKFfOOJz/GR96BvUhfAazkBXeTJWMwFugWsxSTD/RTeaqM/J
dH23fUYR+CO7LM86O7Ks04RIuegc523NbjoMsokOoqJvmPhZMONvSVhBZynT52nauumdE+tndevd
JeyIZ8MGKsS/uIkXi29wo/5Zg25URgT1LhMoWPmJdenwfXaN2PxlGQMlfpUN/cd4dl1BmCfubHz1
CB2euRM4wlJOYvlwxd3G7tIBhLtQGEmidRBWbd6kKbsu0lmEHfYNWBCqsC2vVbRd8LkFbZAbRkRl
eq8V5fWPBvyE1Popv3tJ03Qsjshi7NQOQJZxdmmjgnO0Vutq7JGJ79gAYyImAgDbvDced8o2x2IA
KTSxInxp64bW49OFAIqw0XyJbu8j3qMUXacOMp5uZeyVw4HzAX1atM6kZicaqbjB/S75AypFCBYR
/Lhtlj0pRhaBZ5qtF77dXjDo0r+CfBnhPSzvC0dSjRSkvAKMzAlZ1yfn4H7Csn+6zNmN7Afr3g9x
j33cfbv9BZWcg4x8KFPHNVMX8YXepKsXXLyMJRQLc9/65aykhn9RwGin9ZZyqRt9DM84myk8q9ZG
SlKAeS3WQGZ9VymvRQT9TTCy+FGdiHZ8fJx5BQ61H6X8Z2ALWfBy0nASsVM1SlsilQkqCA0azcxL
wdxa4mxVqlMcsumXMxj4Ls1ANmna7pcAFK2kY9wkW9WaBbZ9zbqJXoLLpt34UHPGPeoUrqpte7Se
D0Np3ogBVUjsuac8SlbOi9e0zqWJ+qwDw9BhfguJzcBBI2W7DpNr9t3bylyUeo3buWPYZy2GbjNX
BfbP2qGfwJKf86gB/pI1lmHtMrZSqJsgVz4jNWG+j1jvSXHU+KIADLgaJUN3I8KvQQ9N65QFQFl7
WKCr+3r2QvahAUi/jYZKNMKgtLZ7IMgL/Gpa4pcFrQ299u6jpG4kSuEipL8ZVznpgrFMHCf7TNRl
+GdTuMjRsQTBN1lAzSQC3y5VCtbA9lKqQChEN8cQ0JgntyKo185TKgX1dsoTrJZlKFVB9yhPBcz2
9+GTu8NMmxeZQwheDSU9b+ndFO6K9BctqFJgEhrnFBU81pmuLSNAj7BamS3f2KQkUdvtjU+GzXBe
CezzXRAL0r9GsD0VJ8U/atabNi1PY7OxUrV5CJR54QpwkeqTeuMcStctbiBm5E7JUWSrhKwV56ae
NN1lX2brHTQZ5tNVUiDXj4IBHBfA9HH383g3NoiM8xPuPkTIDjrYFZApvV0nK/RtsMP2Fi2Kcw3v
cwIlUSfPkLue8DPVBb/vWH7EUtJkc95jB4LQI/K0o1QQDhVHRIB3q5zxvYCihGGB82pZt3gl8bdW
3kv7hJaDTjyaGN4tcSThlTZP845CRGTvSrmfMSzdJqpotfGIbcgLqFlRV0J+AdenPcFX11zz+sAm
fZsq7N51pRCN3uuEJNAZptPNBRE6IbyDnEeUdye1xej8/p6pq/2I0VBFlap8ypfWsgqayXIBNZcr
v3t8ynAYbuOPt+AwXTsvoBQICi6dA+aUY+is3lhOsu/rDgKT0uHWZBNoigoXexOOKwZ2wAz0b7lB
uYXyoQAWpC2wepGFPTVV3J2VHcfMrENOhPDmVSzoy3kgoEyfJfY+F6DRdLkW745onnR+yvyyrNBL
L4rCnjxWt97s4zNR5tcAEK5y+votj2MzsJ2t8utguPJjg3vlkH/qoKQHf4k2P0Wm3ViJggRBzN+D
6tbmDGo12MeJQWWFSchp84Vjdc84YH7YE/QmBpMWpPkrZ29JUMtjibzcFtRzn0JCQponyetGK/K6
KdQWty9WUpgnMygHkOBSwFSckRHjP2ul5IJcsu7KY4iEpl022foXKdN53McMJvlwZXfANRzOqtfE
oEw2iGZIbRxR39jjXCRTWSq70JYumtyNh4Jiq5q3ZBnTkkslCKNANNZBBSm9h68Oyx5WTnfg7VC+
nCrwTf2RE2joaCZ9ruCwP+lolxFjmq8ulNgbK6t/F9z+BTHDHdkS88gmhRTSEjsZeGh/uZXn65Gw
GRDSKFWeR34/CzSDn4Ly4CMwuBN9nSLE9mqbXhuJT2wvO3G2hxquLOyoLiwsvBjhaejsFd3QN8gD
fSvX0Nxrqvl0oA590fx5cKf/+wsLd4ekAofb8fLAb+i6WnuBfmDgULbWRDkLxSqjwBKkMV3eaA4X
tqxki20Bwf7+EvabbQvoJQiqLFl9A+ThSD76zp00PMjXoDbv/d+EDISHtqGmZFOsneDsVi9W5+xx
/QF7Ix2gHwjjCGxpikuISfoq7za/0yXSwPnuIjAH1aFc0EGuT84k8EZ6aINc0bdZdKbFwb5VSpzE
WAV3viYT723BnLZmyK7PpNw9TDqMJRLbq9wAPA2nAK4iZpLMVo2oMrGfpGzu3pTbHu+OiDKtXmNf
aGXiVtnL9W4ij0ke3AHg4ydufZGY4BzUa4fpxzqqhiswIhFns4Nv40CPtJCOqEVlmSSrLNPG1srW
EfgfA6++zygmaBOOyxTGz80HzvVbjqq+ZyvGTfqQOQy3Hg9C7HY7hwZq7JVjyr0gWyzD8lkow0X1
14GcIsllu8eoSz5F65+2nUGv3JakW6ogZzjKsQj7mmuzvmC3tmVzmly1m9Rrieq0kL95yh4/uwh2
rerpimtbKHEqyHWR+4z5XRzdrim0cd7O8FKRPJ8Gk9U2kTl/f74yxG3Cm+TMsWt0a2vIOvfRUZ2W
HK+IsYNlJr6EdwDPtMtYpfaL49jx1HS5zKNucn1tlMVabGR1OvV03ar6IRiAs4BRaLeWb+F9cPCy
Je2QNAhZ4ZtJp1B/9faxVC5pqlCBmrewga2lQ2vQTfJRobssm3kMtBIyYKph1fEKWORXG78Pg6Ha
48IVdd1bfKRVPGYZ2mXMyFC7aft1o6NZhpxWJFVbccWsIoWRQbvxstPfpepwBwAYpjSVeZ1Yp7lp
Jj2K7erRv0FoekK0CUnfcKaiuOpmI9xy9H1C13+EPDKQrnTwOr4bb/yeD0GMNS5KQFrrjk56fx7s
0XRMjjCOJ7dS6d/vEHQQsR9nliFppFb3/ZFhIJaTcKAWWI+gsXdcTFXRoJ/mbDjEN4CfHfOPo/5O
6dt6fHzQ5TfGYHLWBQS07K2mlw/StE8rhLeOQ1FR3AzRcOnWVaerAK6vgHXZHa8ghVd5/1gl3EHi
mukn/xWf1cEo2QzfiQ8jyPyA1Jd3W+XVX0msFVQPu+apqrD1ST+u/J+uWtjCoHHFmFqDt6+zzg+z
YtsW9eWBWiTstrxHpYqWW6utDJSx1y47gtDOpmtRAZ0JCeVEpw/Qd3vNnvjkUUrfmAmcKS3wQLkv
PkFUXKjegMveYW97tmkci3YkSs2SVSdnxfit3cT7xBGhZq4YED5jaO2IUif74lmq/qET+TxGxDwg
1svnq7LPhzU0om37jTlYw4fa4eE+UU2EPBykZsdr/GLmhFddgu5K1ynVbQDiOR4diSBhYeBGGMQg
ccEfHF0IElUlAarUQxJZmxyl6QO7Snj4A/TFj9oeKOPF/SxrLl57uhYjvlllLEHJMKhoQfdRUym8
LCjxUrqAfVxf/g8HoI+Jsl//NufZ1qYy4dB6IgN6ySyim5FjmgK4j4Bn4LrYS3mB3WVeeAW4d2I4
Q9oi6k6N1J6Rdt2ruR6FusobXlnOsQrtHMo/tHfqI2eWmYIAqrVaToJUBEND9YmUvB2Pvys2uLLs
6CBDyRjyGd4QV1i4PPyvTsM63S4Lun+6DoACmnRcdswjJ2HlhddSqpDl/0FAU6FcEX8SPgIJ4c1A
f1BOciGdKKVx4NTVNaVmJq7tSA9qmC45ktxYQfYu+Y3bY72OhDyl8NZCVKKnfBjSwWjCszOFOlDo
D7mDeV0lIoRNDwRl37g4JYsegxIeb8n2QtPNBpA6s9zkMwI/UrWTCaifX0UfJXySAk7gPDvKw8c2
Y1/tfmJXnSWP8hOx/MKqurtUCCTura3nQK6QTWFWHLWrNveIbsLEcs/DyFIWo1HtbDrESLVgg3eH
FdcixYFgeUwpzeEGl2cSbwG600ax7jJTgunkdc3YsrXvsou2yAEFvLp4kpWMpfNFt+motjXgKXia
5JsPuYETn4r/3SS4u2FJm7SSPslKK5FawKBoHv9hD4Q7lAH0+I/pXXmvo1G1FN9x4ETAZcgUWfIt
MynXx03b/FWYHyZNp9xsJbLFIPfTGc4qz+DPj+JUIvcR6WqViNHKKnAiDw6eylVYl/fCnWmIpx9j
RessM+H1zk2OaB4Stvqv0gwBnVeSvTQewo/7swYWjdaUFBQebT9K54sob2uQwGnGVe2BqhIjePMo
hT9WGE/TbPZpbBx1qgR6AfcTFizpqqdXUX/+6MzHOmiek86wmyQdfQlZWCUXh+/AxBW6oBKI7TDg
nJwcCEvdZl9aBRqSVlIzf5MxVKgIsKRTIhO/gf2P+i3aeSdPZ1qbj+WchEvSa9UDUMWYOvuFi5gT
lTJUTOnf7JKv5ISl00+NhCJeaw2l3DMagr6wqpIeE+bm9MvDj+TGd2+vNf/Cze8RLWK3tOFrCCBC
pJDaTxPz2YGWxZ3mRuhVZ3gD3eTnCfq2yc/vtzYjyCZEde1deKit4B1IhgH2j8BXrCJnmUALlrBb
knn97SHHFYGT0nuVHFP7hXKbFb+3Afad7f9XxgF0J1v2qs2Jixwdn+gupEzADYdhVObYC6rJ/FB+
tKwAhEVZjKHZCFvxhXz7XqDhhevpLhEg40OmadB6xFzB3znX1gsMXyoRKTIoSEUTfgIcxQ7GTcP1
t/c+M1lbLeNdeuIEUeqXpSiqjYU+aEXfnXRup1QJ97GMdH9TntEjd9tiVtoFmG6clTpojREUZj5f
KaNNAhmPRJ/Iw+HMG7ZgHWHffjJ7VrvDaSmKSBfgqTp+f+TAtiLl1zWzNqUyEY8p+Cab0Nk/pPH1
m1tSIg/LInepvEZ1xQHKiEl5up7Z2zWSQln2ZJtq83MYU1cyMreLvYa5HmvTqN+k5eXJJCYnPAUT
itXB4Z6RIYgC01ErCrFxwq7UvRFmfYnK+cqq/Ld+N0DCo6s2NB7vtxzfN0FksHyw/VTbpkbb1uJT
vWr0IycF2uipaThtpn4quKRLSa+aWdReP4iskLA7Ub27uAZ9WMUkw+bh6gutvlZdgNHe+auPT0V8
rYvWg+SWAven3N/JhVTtq3LzvlZmTq00woiTKHiu8iGcoUpziRYswbUMyr5VL5/C2kUy+6BGfEtf
At6LMDI9gMXqMNUXXYD7WfkNbqbyDusdGLUue1oh9CVXBoMaU4hH2P6EQcgYoqanYGYWWOeFHJ9h
mAw1lrjkX/QTLQL2Mzlqvz53p53BKUfQoHuab4cVXyygfWOMgJJnMKa3bf3WgDJh9Hu2Bi61ArXk
BYrylT2MrHSFDxCUEIBnMjTwgntU2vMlsHxdbRs/kyka65j65v7NwkBVCS7lpK1EamvnWlbkJq2x
MCtbUNsb+F+TmHx+NPFHbkYRlTTN6N0bR18BvdyGIjLcKIepg2XBPG+s3+9ooyEjJTGzPI9MT1Ov
B/HtpWeDE+Y9oYOIuoZOV7CnCdJY21V8ghXdo2HHmPcbA5N+JyqTmCqKdXksrBkKK4ioBbwDdXCJ
epgElzNZTXb0G/xSkxhV058iwudBlzGUjh7yvCppkqWAbFh4f3vGYTHoJJTSGtUS3LMY+lOevAkN
stwKgtiCplMeR0ywXWRRO7aWZ6sasPPDUxoWtrm9m6Vx2A5y2NBQmvJamC2wLtaXSuafNMgVW9vN
3OnlKxF8cIV/rFzpFWn92FdTuRQGhbhVfNVH1SSDXhDXl9pKs0lyeZON6m8067ZclUnRBntDvkzR
xk6eqjO3gyFdTehYUNtcGCkkr/1YiC8hFKEnVgBRS4d9y60YiZySOjYxm2K2Hsz6Y4lgdoZitWK0
PIeWgBMcCgcvd4pmTbxYplbqUIZLpD7fwMbGEDizpd4iLq30oJS0K4FmwdiNgYZOd7HPf4+FT91C
+f0aHzlIN5VR2XidWrLUDdzFqq6P+albKbHAZ7XJLdvBXVz2P4yEiV5EtFbQne/1AGjj/BMJnpjQ
ABNkoiid50DXhQFwlztaWhllG6jUcOC5SOMhix5ZYehUuulCfjCMSH3UCOEE5Ida1okOw4i87wFf
60xRn9DkkbIYe5gET2EhuSZ2HZIJXwGw1EtyABWAzExpA7SIsCXlv97OdusMIuQHmMr6UGrOw45o
6Vy7yliVV/KoyujP4NtN4Wjvk87HPC33TFVjOJn5jcTwkuCsiyeZ//mF+uNIc2U8nyBaRHgnbxM1
1HfsjhAULc6dxQOBfki89CFVTNB/66bQ0AtizZ+uBT1FjHPLD/qjrFjlcoh18N5tjuKfKIFWQOEO
aIgV21hDVOkN5VZ5BDyeiWJrIwgy35elwxgc3+kAjDIjLRFJgnUiZKsSkWhNFq/wf4Qa8YNq/hnL
2XYDXhBdBXS6Gy3t5gtg1Rdjrc+qo7489O1UPdyPylcW+JPCm4uCVMapJIZb9diJnqjALPqi72Ja
SFT42EiGyDwZMaNbBbory1hIPTLGmUcD3fyqUia558tXhGdquOJE6txrtTSyu6JlgicqlNZXYRe7
Lrj0q4Wxn8TkyIjRzViFKNNLa1MHBihc7COdRO87Ud5JC5iLkaaHszT+O8EhUq0P1im5l6sPjHDO
JFwdP8WJoMmF2cnk0ZuKQCMEaFl/nOYOfkXsPv2oPMqzeMQagpmBqP3tjmcGd5q+UzH1Zryg0LlO
58gID26F2XEvDPLmZeAUAa13y/p2wgDa4yxWJ7IFuTEj+toXqlsigAUClhWNcMhPIecZjiRp61Uo
FLsn4FYxa3oszkXiLvP3MuglRuTcTB+vKY0hD8GPdntTW3Agx/EgBNzI8Gt5QACfJcnUdV/Bw0aV
4SvUxYSKag3g+wLF6eOfE1/paB71EXMA636gWUVeR1WBTj0kDaNJLzdWCWri8YxVtRKewTyxjLW0
rPR2GZ3V6J+SI8eF0lw9xnYUxSvpb6BTESyROxllxA8jMSWbdChU5g0nK7THApsVB5HGxs9PrhXJ
DboUvWvKlAhh0s9nTdm7rTHnBX+iwswtU6jewbXQaSVQrNUL5K2ueUxgnBydOq47h72aCMNKM4eW
7k0t2xlcqp/ejlETdxcUC9KgJjOa3Gzz98ycDN8dNkB8GhWtOy5dAi32/jeHtUP6PpBXRynvShSX
OdcRBzSZTIkECFxDCpUYiTebmO20oxWac/LFfMspKbZ40DVgUjsinQPe1IYWB/ydWohVP/n/NaD8
laM4mynE1Qsvtp4o2+C4HPjf+qNClKc2vV6kW0h5PIf7HDOaDWah3PbXsbO6NqgU3RyuJEUXSNco
z71hN7/Mtrot8Z6lhAf4DxiNCHCCVw2tkN0IqbSuuvxr2crkqeybIeKWO+Pc3WyQmHxaE4fl7CJx
5ZS6wRR8haQYs7cA2UOHZY6/hWApMdB9jtemd4DryAbbrQNhU+MH5T/NX/u8WkHEuwYmgjzYIQJ/
e9X1pgYxrX0Wjdcz/G3iF79vjcTu6XNyK9tRCwwabjEPJk/pDCOu8vy7X/NghtgoWHuH5HXjFEfo
iZJZ0p77sGsnehLepIIvCdfSS6jsa/tUd7pyTHtcEzcjb9tdiAzBBdRX74yVViwCh9TSgXO0CyC3
NoGKaW0Il+QT76ZLnUrIuAn9yVZCPK4Ob6e0aPO23JYooF6ELKOz/rAcR5XPgvltONesH04xWsDc
ZOvi9aodl5gJx5W78FJdd6Ylb4B71O+VGhmZrmr9ISmvIdruFXOqS2xfnT1wwHstyRygS+sVPL3j
qJMWe7KxSjoLZIdrVhaR/12+tMWEfHjkpNLFy2FlssJUsTDhbYJQDUhFKvaXW/Z5ilzmZryl1XbE
hVnhadTmOuyMmENpB46Nl3cseYrbKsqi1+sscXJCIla11y/47fZzDIGhnY6KV6JLHbG85Y+Kgtjk
QjT/F97M+sLVrVZr30PUTzGGM21IAMPdzPoBd+EwnhokCBq2Ik+AKkK8HdGeGciUFjody4MkTdDU
5/q7mokR33F7YyVg+HJigQ03ajxZNGDpE4J31N3yQ8Ob+yJ3eSlwURYA2yCQDb4tjYyVzf83Wpge
B1fQAGsIV2/dVjxeHxBYd6pDFHsiS25SH+jLYkPEeOinsZcDZ+0XIYBlojBU3p52qESlDrRAEEus
GJfuI3x7TPovpYZKtBnYnDXGNKYSbXPCP/1dVURGbjCT48JNf60wPeiUNZzPQbGqfuqAdP0c1YPK
LroCF7HHzj00GMsv7aEQPjG0+3K3ma1hKTUgxL/HOlwdbeKZwR1B4cj+y8ptYHlfku4isTdfZNXB
zlf/CZkDnpJHrjwqQXtsOPR6+mf/r8W2LUm+x/vYvMq5g2vUNUJG347qRnA59BcRW9V+FrlbLfNk
pDPv4bNRsxG0Air0g7GCUToDN/VGIytUcnWFE1kwCLKhL11SGCfnv5QOEMzYdvPEXPaPQ11x9MJF
xNhBEvbsEBumdke/SVDrZ+yRzt7eug4tPgrKZP7FYf+slvsl03kY2+7rcgK9aNQkzXExtUc1THHc
KCVNgAvbFW48azai0rVihEOb1/qliaDzfKMz0FPkL57T4muo3JTow8q/Rmbg/iRxPi7/12XPi468
FtaIvsue3q0Kb6po5G1gZEEEj9/38pp431gQG7C6vyWR6oOyLgdDNcJv4AGRlgUWYp2IOejUzhsK
9QzBPi3pTuDIEvzZaTVqZk5t11AQfdGofZ8Ugg9xKR2vmEqXwOMo5EcaHRrpJEdJyKd7NTza3lWP
OLVhO+NqgQBtZjOvBu5HuIwGhn49CfP4BmK7xiwxkpSN8Gg9eP+TmiBXWKJbgybjszF6A5/aUeYK
vW5Vhh83XRoRsaE72Wu7INdmnc3ONu453eos4+NwE8BT8AZDE4gCbwfdMtnJjWF28HpNByGwmGYf
QVF5LkfOOuRelE/3IVBvPG8PpSEucmSqc99zuawd5iL37DhdDaesOG+KmYIB3spxwYYsDOBr6rXF
6EJq9VBUVu8A2rR0g73t1pFFRg+9nEFnCTjmuZROxPRn4nwmYSeZBdEfC1ypb+EyFyjapHwk4816
6TygYR7oMS12kbzp/oxicp6sOr5NflylLSCI74G8y0lGBf2u0BQ1iVKhAgRl0/637Fs4RfLIrHdW
9NgtfQ1tw9iaQebHEzLB3rWJSL0w6vMy1x2AXJxOQe70DMIDo0gfh25bzi0esTl37yb0arhcovCT
b+SsRpYAa97zvMC0+haSnmjJNuTyazdsKotZNnQ/iTIiJ4ExkKSYzf3lGG1KO2chBGLSrPiJJsuU
+UU+J/nyOxAxVn6DuQouvIlLZMHGfzG5cAM4oALh5Xibyr6pZN5BheE49RwpQmMstILSH5YDnJQ2
/t0dp6kNtcfsIAw/66V8PvrHCAEMDosrxQFRJ79gTY3CaVXuwW4SA0OCCGbbvXyzdVZdLIbRDKsc
CUz5aMrdlz6aprO3/8WJjLOsVANnlZW3Oksw/f0AcOHKV5NysGclopU9cdpOftwwvO0SgbPqiRGn
8OTC1M2Rh7dlrebaMGF8ZSiEs7DZaESERXg5bsszpenxEk53l4X6rqLXzU+0jDIEGX/XvdRd4yAj
kfwBWgf1B1mBTeDOVBsm1jlAnh0JyS8ppxX0kzwnuBZV/0JLTe0f1UwDZruU6j0xEfbacbqXGKIM
9wTXrIbzSsjx2sjH9ro6zDPqN7sp5grILzJk2jNsYqUaVrrAtmb+oQoV3K0igXQWoZVaGdVOqXYX
+59RyjawpAw82peCRCkGSK9jxovhq6fdtZniPZhRET7hC3OCd7p+tQo2+VIQq7a3Gt6ku83foivV
Q6WQSGxefLKt2DWEws2VIQGva+8l8XLt897JW7yBrrwhrwSY84aLZgF/fqHfRM9sbLQ7Xqro2D9d
AohhpnprenEbiqjUUqW/6J3MQH8FEP09PZf5h7i/vjLTskqrPN5876I3ATjnDHMxaxgC4ei4vZsn
mtHX9RGkmE4EIigEUCfMqz81c1b+JlYrdgnXkTCKzmN0W2KJiAkmHIgSY4LleMMMh3ZdrgR914a5
WAQBNdwlqt0ywcOMaV5s4ifks25BjF1TDMasQztD0JedC89ijqGJ/Vu13/XsL1BA3uR6fZdzg71e
0fU1bSA1o2Pym2griKGLgt0HPD1RDsmaYzksUeM8Sj998afhdNQwTy0WKSyam3+JGFtKxZ4j559D
Li6/l4GupGRRBQ83iZly5af8EF0N0NPloa7IqUcDWqY4xemlcyYK0TetEYY15nhd+weu9ZjF5vZ8
2NC86EwTjupVVrk6Z7xIFxptfQloo54lVK2w41fE7/p5QEqY0aoyoAcHy9WQYAIzAxGiJWhlsWPN
XBMGOVUqWl5voJGfx5i9wSTq+0N6gy3vJiKkiZCJVU4jLjwGaeEI6THAp3ByuWhHZ64DAP4FcrzM
l4GidQVZGCRPJUM6fCh+E77CpmKRZsd9x4VvtMj6wZR8HnBMDdVnSfXgnTIy65sv0uCIXbNPxDT7
sjtfBBTsvJCyO6KphQCy7ZumWDMj/ORlc/ZvjbLdEJMjBvUAVa14bKOvSmqF1j+02W4IGhWYQx5R
YdhGiJjdqQM8NLTKU2Srz6o4ucuQx4k9Pz5zZC5Tq/odgw0MZU3xMffbK9h9jG1XVrOlSsuK9lnV
CyZfhGeNgiOIOM+CCshcSq2t8dsh/cROBTmDYtTCDBUe6hcqN30RzshljFOvIQISq5iFdmAUhEMt
DYbSh0bRYY6jn0u5OBt0qppa14XgsOcgGNyhAnzQVljitIBCzAo0cktv7Ua3lxWAVQGETMvMdE71
uXHhOxKWlPXGfBBzCBGwEzWvir72C+FHfnfmXpwDXyBaxUP8+DrFB2+RVbCtQ0/BxiHmQFWIlNhu
go46gmBijtvTE6sxmEf3AYERNLRu4VJocyVPY31SfEFLzQnHLgIf+gr2bCNreXJUCWbM7JLRtvpE
AQytUMnK3n078OtAv3mKW6xyGlPXL2isX16nHl+Zx+f13mMtbo8PfrqHn4r46ujFgWaMnivVi2Z8
pjRdOa/mAI2xJJIjAXr3B1bjq8DFz66bfMKHGC/O9yHwVC5U2hHPH0H8zLyckVUvxkaOddGD5O/Q
wneq1YMA5uN/KibgFdSjua8lZiyg3YpaIpyedIo/JJwdHrHVmHfl8itXFu/QsuA1mfI/tvht3jBw
5TKyjV6DJOXX7JQm+knMLLbFDN+EXGmHdAaYAHpzrm0T3d8uZQYgA1Ctz/O5FcJb4raioL0j1jOL
k3ywpqhQedEbE7sSIBaCtYpqY0QR1OS8w8CBVCiDnRdZIdNllfSTUfGgn+D1CG21A9oe5Kt9SGYP
4lUGmOTj+gUol7cXShReXosFEVY0YP89SRz9UuAjdnMoMle8fKpRhzmJ2ZUAIewYKOkvJlHKaQA/
p2HbISFBsLusPLyNreoCQgnXAhfRr/ptyphVxHuz7AlKw3fWi04XfYngolVbMOe0Am9NnSu0WGCQ
kudLRshinOts47qSC7SWATwJ7vVXBB7WYdCRbaJMKW964nyg1RjMCWAGvKYmVDElUxN9lbzP3cSI
6HzApWhCYwSoQ5C7U+AdoAwF3gmbtDIm7HPYMRbcnb68iL+2bPBS0/Q8d5uIyRQmPTs5gBh4MAM4
ay8C/XKs1j7BGHHfc7RlNzOKY3q3n7Yjle6ZfxDth7BO5eGmtWj5BcQ/QTC45RUaIEwSeBBgh+qo
yX6+U8hl9by3j6X+Wr3+Zk7upmy7bz/KmiN06QOHYZ3KDrMJ1IHYs2DGgZ4QwPH6l1Pf0dbITCKl
iDVW8qqh9jQ8gpmmdPo+rL1PI6NKYkGzqORuM/D+mzRA5ut7YlaT0CHlr5siD8bAyowRv2O/fMWA
gh8j/B7NDN9/vJVGQrAfUKorqAX3fL4Zjc/2HVEePyFx+StbSPf1brWurhOXqbUVe7LwvL3JSBJX
gqbOcYCaqe9/VTJCYsxaTfQGFliNKPxXSzqWoorr1vJM5q59hDHJK4b1SjN8eWapOaOp0vGQNQsS
qOB7e3YObpeCncuAEmWjV1h2+Kzn6DO35r5TPCqV8DMT7/hqVtqtnC9uqf7Yn801hEu7mgOqyFqr
p1CW/AE1SB79wOZ7zGiFeemxgALGjUF0hjQzLUCY+UeVwzcsai6vT67pRJY5i1UOrjvUt2D10DdO
juu68XQH923oMd/JunUp6ARJhey+/j5DbQD0FLANu85z/dEISiWCEW2qFM3tXYBDLwG1tOiUNYjr
MREhFUodyBZ0cWokVALM2pf/pSoMMjFJ96LchHSS/tksmJ8hjHU1CUP4ZLd8Jz5v3d8b0M+Twh7Q
mF4O+y2NX5gqQBkj+Fqt+dY8vdG4TwnnQIKKaYPfNaGpiMWlURYokQP1A4DnFk2iC+MDuYBFZkbv
8LmU8qwaSwXHF0HDkUdFdQVkgthgSE3xDE9/SOkH3LMrUCoTvfBJNvMBzWdq79QFD1dBHY+zsRnd
5yr/YD433wMkSd52ZKuJVDf4f+FTmcY1PS0EMDrBRSfAhrn76o5Z18+mzQS8+sMRGnT1eoDb4JhK
AOhsNhLIaO8ysCUbJIHr5esZJTa08OczwCRvtqxJWfzwlRCGH+Uc5Pt3yTzz5A19LlWICIrMLPj8
EwtAV/be06y180lM1G+TyuzzvkQFDEpn3YdaWmx/hfHmRhlBVIZX0scIV+OdRVl9Hx+9nmv1c9NI
gKy66SxB442yS1bw7AJwR5Qn25i7OoBZR1bkybSAyiHOOwL6n24Oj6xXm7WRab5+B+0gmQvrKn4l
KcfhPYgzAjVwhRdQ99XBsYvktdxr2CMNzvB5Nvmft+UHLhQQL51t59sxwt8lYYIBO9GqxuAYjuzU
AaNdSY7dnAt4f012eVKpIdrbBF5geXrxY/pCRm1J0SegpkKrKUP3vHoyoHePs1Mau6LvCXUqq8wi
clbj3n2tOLBwzA1rojeHKTHeox0rSeZ6VU1kHSQ56TF00ADexFZ9T4nbTa00kjw2XEKi3sQnSfOk
01NY6CnqypGraUf5nk5e48ki05caCw2qrw1XspsmkwPyV2o4LIXGG9TVvNfWYZySfs3WlQdfZ7P3
1TRf3WitmrGYGD2L6Tu6HtVAljGlFvkuI+lHAUdEGlJrDh1U97H7F5dC2NA+KVsysd+LJ4RgnjwF
0zpp5I4LDsMD8VyVCzrNRQYpvOO26+TIQprbP/cR1MR4alwI7DCZ0G65Vn79lggvM7AfYCqsmcXq
G8OEcBsFAvIsHCbywDaQligZSeR/Ok7yIbvBHmsv94eYlR+VgwqG7DMrHpqxyLpoXrgAZn7UeqE9
TtMX0IyIjcdrxqNNdP+U9K6qps94zjXmWfoSsYEnyfvSBsbcJn82WZb83MWqECdi2WK1VK40G9Vb
9vdB0OBxZsoO7jna6mj9jZukX+Ml83G4uXUhefD2zkvTFTNQ5H+kD7QHScQpUOaX3M6LQ5SnBrt+
fJ4an4qr0rv8Suw9T1I9WD6Kfpe6bBPOqjuOb+mh+tX4Rt16MPqcNcF/f4Rlnz7wN/fV4ESoVfFl
+FCPT4i9ogUZJUxEbQaih5pLAZEzm3tPXBZSlY1l/CbEexjRz68d7mqcm4Yd7NGIl3ImUcXOJv05
ATDAaUwq1181VAepxJHfLivhcl/mmUvscU8G5kYiPsDJ2ZejernhIZux9W9PIbgwa52NyKJpNIKh
iLsNUFcCqCr1uF9XXOevl2FEO83PfC9Rnjnh7cjUuLjWYjpgMgzc6m0aYwpHc4N1akQHvO+dfluF
L02e+LwMWOvDacmfoLqKDsVTcqxOqq7Zbl35kFAgpjY0/hcH3UCidJ8gLVjzIIMCOEKS1fZPIekY
qBXl7l42DYHY+eJeP300gUmKaBFtagQkvL7zfkIpuGvodU82Ueu80B+bcXITHkcXHwsW7ze3O1XA
RyGxeP1VLbSncpfQwo6NDoEEe7JFDBjBletCDRCu6E2BoKsUq/dgVM/VZ16Hl8VKVXqc3jt8LmlY
v9BZNOq91amdPMtjxYik12Y4Sr8O+ysssi+xAoMuiYW2VxgEt4og83b2rqfKDzyl3lqron/NGrT3
AP9fF8UpQb1f68DgRgtTI9s8p7n6HNa4+aB/KTq547RwUY6rAAeVCrPHsvQJRshKuzk00Y60RYpZ
SRu8ln02weqCgE3iyrptTiRKJZYJIkqlpfsNVtNZZxBeGdpDdwBZ09W6v4VjVK7uiB6rcGYf19OD
+Hx6FXkFmYVJDqgJbE4826yN+A1FWVOQGpxiNPQ9IFcOQ7zEP8eHtJ8RDZkzywYW4yRBuNyJdYiR
WHLBLMeh+yp9T2WvYUm0vQw70pzJrdeWijWERh8dQtIVREiN2s65FBiWyA6TgIZJ8orkJXKEvDl9
m29tPuokZ8IcIAoDUYQIyzZLoY6ORVklZyMo9mDAmIJOmILzn++09BwczQj+y9EoviB03Un2ASmM
zHyFYaHQmmAjZ3DBvxSOKNb5SeqbT6TGtZhcYw9RVWkMHn806QdLAbjMPg+imc0zYgcSXi66XCh9
YgsXQS1nVtozcsMw6mZQ1hLdKHTAr3tH/lOZnGEFdYdWBSPCJicsFK3o4ICbWFiq8NhPfS+5UiEu
vHxlc+QhHS+gAJ/yx1YzY+Mkp8M++0exNZXkDTWyjnR+MMSqF9hmWdDUOJ6v2alH2P18RpfUwSW9
m53JcVn+i1KJ+FayR9Sc22efWjx72hSF+ydIiarhcGum08RJ222brsUbva57fpB6qgniSVzYpvKx
BJdeDdWyaOyAPMsXQAOHzXR10f1c3v+ZbeJ/5tEzARVQPmys9jC5madGRmSjOVenX8ZJWqiKxMLv
RRA900xorSLVOttFxbB9zf3xxFMTa1X3i8rLgaR6tg7dHaqJi0RXrkunXxYdGQJzOoTYSTb+lXuO
88OQwo2KqqpoZ4ddPw/grJt6sisimtBsYkGySwjGteNia212DYC2bjaR0b+u0UA3FzhOnkkJLICN
mKeTynZdOzd/2AYhBOS9uxB7f8puSosSth4MH+p1PySZKFUmcdZ/qRf/TpHhyEsLmAJZwBoJkG+S
6kLE+3UzmdOmMpQ/IsVoXgJuzY6BOwc/1a/Z00OGYixWw9ngusEQ6LTCr/7rEVK0KvHpLKHwsXks
hfZWT7EBF2K+9Ti2NkMGbhMBQeleA1xHslHeqGQkrcIlROHfdu9imA7qFOqJdFm0uO/5drGuj1qH
QBufI0qB1810prZAlEIZNrhzijo7KouXdw78KS5G0KBf4kP5CKE1wNZZ1QWQDqF1j4PW2nMXRya0
HLApkmaeu3tyj30w5QEb1Anhx4xL4s4pIRd8/L7G5cvQZ9pWtX2TVLn60Tc9EvtHqzvL4jt2iLi1
BJfGSdmXfdQcOX1rWskKGpkMNlElObZ4jK9TB0jJLCsLzyMmEvndgMAx60RnqpfPUoLfDk2h3FJ6
bEKfGN0hJpaSdQ+VEM087ekFjSiIAOM+bvZhvXX0UmkuNE4OF79eYZXojBIZ0f/FJwAUvUh9fbLc
Xfr/4tUKrcoOfldznSsAIK9czSz3LJ69WUhxxvdljM/q/kpM4CgajHBWwgPnkmPuiC0O3kLkGdTt
nyISAhIjw85UNZyxHWK4iIuhHlw9RapEHG5bYlhECkuyohrR5NS+SVrWgDPPPozOtDAYcAZrlNC7
1lyXsEM6Tqtjsw1Jfkr54r1KM8ghY9yFuYFJe7jSLjPbdZKTv5rJF7ICaMPdaj9sr9yszXW568rA
OZSQHU8MFoJPAIJs++YL6vnrF8/HlwEZ57RwvkKbwb0q3YaA3mnABSI1em8BDVQClo5IyaIiduvM
AJpvrbd+uFP+Hwaq0x96u0xVsuJRUizGhBEZJh+XN/Vyp4gjADU3NKS0d6rVki+3PT7fN+nBfQjc
J67MkJjQ4a0Ca3ycfe8DsG0BCH2oGhxvoNyvfVPRPbkaYQq1P/UWAAbJT7bHl1195928bQauD2C7
U7yNY2j2OT2SL7gmmaYypQGGpoy1IBKYYTxFp1NcmiQyRANoh1i9iQqE0ZxpZFdw6hpqfVxAMNEY
v6wxA8yygMsQc+nlYh7K4FY0OLnBiDYyk9h1HtN49OQEJTKeu+ZqbbXnIGoiqHmpV7TN023J2QyK
6Xm78xwMH/sZK5nFMc8amrihLtD/HB/qBlFjXojD3eOnrCsKBBtW4ilOCwtwkBeY2mS+lDKmg7Rv
4Ne2Y2NeYczOdAWMqQ7w/RytibLcquTnnPogCZdBGpIdh2T+Kd3TatJ5aZ2se8+MJYbAX1fzc1d1
yTFW8eFGPv7hAxsCvkbMZ3udGzqpG46+MS+00Yfy8FY8tS5lMnPGLxQwCrlMk4jFGCFSF6fKm9c4
6ORMyrAXqkg4s4aYI84J9IUdurED53eIbNA/0Z1JlYCAgkYDQzBGgUP6IGyjgfEoBhQGvKPPD5vD
5NNMFEMAoRGDoqRIr0+U2NX6aB2q2T/YKwJbrS9Glc0xDIabAXorcIYgsyK6PHaM/LRgopnDRDbJ
Yx4aM2imS3juRliuts+Ct8vOA0mAYJxzCZNMdYhlrYNPSRSKHe8xIlPf2uJPS/nN8BndrAxSXgTr
UqIxvDH/YL9xQ1uanQUesPrMSYF7cYBT0Cmcr4lwX0FUotvHGac0+qLyOXtPaR6wFlNeenfAACxw
D6xAIMRbIv09yYcA7VaSYqanifviWRhCGf30fNRveJVkM8bRjCxB4yziJ6nrXkr8nROVEPI1hZmH
bI60ZzBM7Elv1JATk37WBx2nt69MKI2JwuzJVzIU9c+yoQpv4Dm1ImH8Z0kpM+dE5/bc+iyeJi36
kIshRsNKabejXQvhJTHSQnh76OsUS25lG7VtbtpKwAAT6hGPj3gknoRYLT6ADdy7G9WitrgSO7PM
vylgM4xDOtHRyZBGzDUh9k3YpzBQSZfB6bfhB3JTAgrB8NWxJh8W6F/UjbZaaAQOhQTfPcpnNflo
bFrZ1mQQQ+JUn2sGkNC/yik1Drm9iaT7yrlHwN4M4YSWj+XMS9DP+G04KNqocYt5asiDIv7vWnNv
OrgVjjSYtRXZ5+rLp2/q1Dejgx/GWhDNAo1eGqfcLxy0Csq+pIq7REFZxpKXaMLenuntnKkoEN/K
fcNxXan/MrJptZfBPm4x3xkbYaxovwYQRZbn/BjgT4l0ppkAGvRBKepyF4BieEtF1aXACPp/wJi/
gJKOgpCCk3tI4c8/9Tb+QghTpG0Dmfcp7P5jHU6U64jQXBRjHKSHR3xMK2xrR1fU/cxCYK93b8Go
CwaYHPgVbMObSa9o16MqyZe4fSMjyEBYbcOrYeMPhsOn0kymTQu3run8QGzGWkWPxlREUAnDkuyF
z4xIa5TTtfClfcKNIs9lxDwgChLna28hY7IB+hHfLZ+0GKZ7Zu33mS13q3xx9Zb7Zdao3GLkY+Ij
k8+TvaRQMHwIm8NenPUXy7SVbWm4qxcnp+BTp0nMTntrwhS5cUA48f/XYSPRhRUb9SesA8ehdYoH
LHDEEzfVmlX3hEW/kXrPb7pVR/EMJ8ll8AGdsRi13T34aAAc1xupLw+pSjyPnUP+aTA05uk9AzYo
9W40mNGxyI7Rbme+3PN66/Fha2KDTsbCcHmG9XaxQ2U+miHlZtxm85Y2vVRQ70HpXpHynYl3jdaz
Xsm77hUuDx0bN619LRAzXowFDniTbv3GfZUE3VWnP/VF0OaJRjATBhyF7c8KZLUpDEhOo+iXb8hG
gIi76UkJRZuhfMgacHjKoAsQdtc8iNYisz5KrSSmnWEeE3d16VXr/ch7iq3w2xihN0J553ShLZ1J
tMXNCrFuAZuUmXJ0WY9H41ewzOJ27u9ApAVP7eiV2GyMroeSuyRTo20UBUFDcjMPpGE4vil4xIZN
HatS2q/So5pRULYJ+JjwZ2uAbrrm91CgJ4XBfDfz7ckWHaE9cgGZkuXHSdo7ZRNvaelDgsBMV8ip
cT4OV93FecdhEq84ttYzoGtl9d/FHzsA+WK0FiqSEl2HhGpHMZzAbndI+cnot3c7pSePJbz74Zaf
CkVwszcor6nwFPoyIuuODvgqpAaMUR2ghHMNakAxb0wCJ2l9Lr+R0WHsFftmBC5KfSNkKszDPGXo
r6M7FHlYG48//X4UjMeSFp9lP3O6CP51GBsiqM/xf5cG5Apl9e+jvMPeit2HEFIlTIAdYRHjYoDF
N+3mJ9tQnFWhlMAgntaBfnqY1THyTGr6HKm9TYjb5fyt1xQgOVZRkgKbzNkQKYXlhlLDtMWa+jDu
ecSzBaJGzwCGiPOn4Q1Pa+iGEGVpaoVdQ3qNtewa7nvfSFL6TjpliBTyYK3KGe1zB4aNeutUW2Pt
14GCghQYOO91VPCpQhZo+jyXYMXt4hO524UX5N7d4fx1sP8SM4gjQwf8w69I1zm6Uuu/OH6gJupO
4KbywniNh4dBeu0oBR/0dMmSF04VEJZmioT2BjsG8aaKZUqHlHwZJXY+q/Z+P9vtdUPsT/ocq+BL
N+spzKkUey3IH4n2vGPnSj6/a5BpWIC5akA38RnsB1/lWSB1UoHjE/c19prUA+UMOdhXHqrveqVU
s05SJ/hEkqqjKkhwvtgnW9HUA39OFxkCAQ0/druJBkCBUNnfb8MYdK1RH47oit6g1DWBCQVfzb5R
cSHsVOljgmzKebo2b6AfhmaUs85KpnGGv9LRnCVIR3KNI1SWyxiSsi0g4xk/DsmLXPbNaxGcHegY
1UUmN+KB5/BcMer/nr9XYwHF9WAMO7TDZPWDr+qopsiHkjcSsc3dhNunohjuLE4fHScKfs2f4AA4
ty3hIePBkBMW0UzCdF8O1v1Z4j4jFPgFNdXqd9po6KVklFZ8Cvg4fDrpReujyK9g/pSiaoQXp0K7
Tf3AsoEJ9g3UJ3ESRPictm1VmnTOsHoIJerZDDk+oDSCpS5h7d3s2GWWQmnHGPDQJDWiFaE9U0Pk
hjjtjq0qadRBh7UR+iFNdYu4Ii5Fw0eZ7gMF6aYhw87LihQfyWhKOjm4tRJfm3LMNyN0XuedPK4Y
vV5m0kKU3YFXnFp0r/oHpEQwda/tAiiY9tdan1bal7k3gzMpZ/MaS6G6qik0QPgRg0OF4BfIDwQt
hZ/Aw6XeiJ4jlYDSoHsV7kYg787mUSEV3t2Epg3tzzTNdzaHkUIQdXh2DNc9S7CkckkSYhx55nEx
VgaYe0H6f4rloHVlcSdyumow9kjrj4hgwxWGCGhyBqBntU+ZqvpdmLO3dMrOLRyK/aZZnU7a9Z81
E+/A4Mr6fEsRivt9LWhaNMv1x2cFeaTxhxSkb/7EOIEzUaG3jBIcz+QpaUybTVSwcwgjEdPU8fZp
S7Dmwvbq04VRlN+AjposkxwgEwwy63UVZ6G7lDXRsmxc+IpcsI/4gMRaLtrk0jix4YbN4gaNHQLw
BL+Vpjr5uiNavH3I5WyXi8cYelexDeopxBILPKDc0KzuiiCbLYtLOpRs4k1I5vQLAS8ppMeIH8Fd
eavkA644fPqBO0Oy7DJccymG88fb1xKQWNWhhc9tyw3HQrZkYcpT8BpjAtN+qxfCNsHBRJ4+WSUL
oyt1SOJcYkq25/QOOrNH0PD0wB9Jjd5YMCYX2jfxVs26qtb0yx+9x6IWcb1GIMMwyhliG7lHoTsS
9zodnDRzm+YDVwcCN8Ym2hJMRtPDWgVHS0vhzbZSpv/Q4QtN7Jq5hEbmpHYysr9H4Zx/2DjZUX0f
n3kVt830A5pUZIsVVxcfN5NZPzlFEeo2Dc1pQlp2cj5n+rTb6bldO9d0kGznPm/VAqPqEOawMT/9
2reZyWgCIqxA/rz9pdSEyWPiQW8xOhDgXBvenceoKGxNLhkRJeHuR2kC0+HQofpVZq2IPgw+7cbQ
9etbzrC1BkkXMD7lfA6oWJ7R5NHeuNuK2zrCyuYySrHAfvcsdm3WJtju5goCRkrnYirPuNEaQvzB
TOiTSeao04tn4M6THj6rQybjRhzsbOGQzmvXDr8TdkFaGYSsnUk7ISaIAWiuRgSwAqgn+IV06stJ
scPidz4P1LJ7MB1JmCRVPna2Oh59SLPm7+EU1S1YqAGBea5y22yQHqooIB0KMeE9qQrbO21bE1A/
bXYT58ehP0ENYFvLATWiT4Qq/OLSKONsymkVS+S6OOpqF+TXZijfGEyFeOxClVd3Jbk6vHBgjchu
44FmC1BBlK36nRnJyefnnrKyE/V9v91CuBWIURv3zqUnXaYuPA8PnfdQvXC+tB6Dv7miilE9Bhwl
OPjUXCoVYtkxZ038BtmOyG1uhEwrzhbJtvfjsvvONEg2rHIA1vIiJTIKjSb1YuaAydbfJj53ih/P
APJ/QVLzC40gI7FXNNcBaUZ5/RCgZLDgu8JX42lxuhSHI1k0yguwZdC9Ni+bSzakKkqpuLJ5uRe4
nGKeRuCDeOrV6tXEr7IamMrPl8Q6pukBCBzsEG/hE+4dmm6N1tcmVQ1nu2vpRXsqJ3kSYx500Hl/
nYfWnEV051hhjtOR6aUbQaF9MoiduS+VOdv9m7H0G1b7UhbQlk79whyikB+yN/TKYIZavFzBaF96
dYYlr0v1CvCXf48vbIw+3B9rB4ZnSMG7H0qu9+Jej+vvnnsS+evGaE1qAljSr3070IZDtFAd1Qlr
ueomY6psIPI1arvrKX5seo0qZOfyqb5glHXTZdhNg/zFPohLWbt6Xqw+CeuWvQLM3HSTPoJruREt
24oz9z7EIYGvdwSCqP7gUHsE1taDIMZiv6DJ5HLatG7EQIKzcPfjc1fcJPCcDNuQiOy4FTm2cT9j
OLaiC2xuoem8m+2HjjqcIgE5vDM+2gp7ridpY7FZvJXskmjJBCvKMnq7iNIxKqEyQ9XOTfiRDlen
1ENAOBpOdb18mmE6zhBjiLifR3x+fkDni3EDwQ9m+apdRXaVj+poZGaxFDa2jFnBxZqdRSF/0hdH
G92kiL9NyOpdocONp/KzQlpViP/sV16/l+U4slDN3mEyASSaP2gQ93onGKSpiTfzyk6P5u3YPr7r
jiAOBGlwaqANQIFLsKThmNWqcm6sL3KjUv+JpdfoXmnSX6i3uzRayu/gKm9EeCXZKB3y+XEYC11p
woc26C7DhKQaXbS/1z1SBiDefk+g+O9PdrVjLEVwvDz9wvESACi2cP8aFPr0IRlA54qP4Vny1Rio
P7tSDOD9OCEzIsiqruIkITcqploSI7gsdGP5iXXKh73JJQ+n6XJXrs0SjRhG3lBE6t82VtgLxRPa
q3bayJqwJFeUeDFsJGpxVUEi5N9wmgNo61h4RFwLLmMjGZrc+KZTnHt0bns9UG6OahJWr/krgLfb
sACBDmY2rjuHadYPgHcd7sBnOO9KMjoHsr0If5i5bTG9eN6OVmami8TSshv/ewx0JnhnFte3EO6S
N8s475x6ISnu5sJRRW0KQuNzvgMDXZ7j+sPjYJQMLtUllxDYCWxCdxF8jgkN5dzA8uFw7VLa94Rr
gECvk8m+bEUmwqMSDnN9GzsCQvFCKZfEpGyYoekBa7GuwU2VbQCfV0T62GvWXW+Y+S/8HXgSFl6t
liMIQigKyB0uo7wIgYb+JZVsNv2MLPsJfVB64DgbTUKgkMPDnbFsGECL5K4tqotPR+So2e8c2c9N
NFMhKhJuPVYC9VC9MmQd3Isq9luuBxLJr2/QV1Myn5ANcDrVGgt0NYBcsVUrxD71jkhU+8A9Yg1n
kej0fJF+C3FTKxYeh8Mpdpgdryu6F0XPyrGe/3Xa0RgNNYVDehjSkhru5NBna0weOIwC8I+W8S8M
8G2nyLIvqxsRZQpOSlXf3zqnm4KSxtizo7v8JDaodYU2hcHDunDa066TU1zk8uSFSTDh3+Y393/J
DFt8Jb+9g/kBnRXnb+XVg3oJjydTldFtd1xL6h2X5cmx9ILKxpGwZ0L+AA2XXBEV2oyjdwOE0YKi
Mi1nZv1AibQIFlybgwKdhdVvzt2rHefO3vDr0oAPtaAffpdxQKObXewuqipJ8/b+7kmuBYcg5Vt2
EOWG8RK2xPA8YZ9mQ6iX3sfoJJxERerTvbU6U1CweRhQtgbhqjpyfJ/MVXBy5uJjyCa6mXJvTD55
F8gjSEGq4nSyhyoDheLDcyml6hMTcbZbhkMY+4gM109N9AkeCg2UsNqJqRO8iT/TqJ5bT22q0CiV
403OSF7nDmzCdzWkRjA61keoqC9aXPHl9mgY61WEJy8xAVkps/t5NBYE3G6PUZYvXV/pcMKxKLd9
6iIj9UkeU2F7bhnOD/Pu46i7YTXokhqlQYQZ+oDFkjrwEpmXWMSDMym4CkYuomufDYceGtdc47In
vMrnPYyFLC3Ku4hsKJPnAWnYMR1+Nf2DKqmlTfF4EtV5mnbR+ZpkZ5zxziW+v8NA7e+raHc2zIQE
QITuMmsFPTNv3cshUQPfIsJLBuZEmQCtFMU4MIIFUDqjc8PlmMubU586uRPiaPme0l+cesvwL+py
QmYjMBO1NTDLKLg7KzpYiWhB6E08IhZuWcmL7dPPPdBzCnkoXQzmfaIe/igS1G1Td4ZpnTLafryU
4OAWdIdbD9p2A9ilMUuJW4aiab6CGjAIZ1HEVSISlErCBQSCm65NkPiz8NefmCG0faxdNuofx/iT
oGnkW7pT97gxBUQ8tClO3GE1s3ayzoDW8VSg5IajezPSWJnqYHcRJx5C8OonhvUxRw1luqaopik4
tmdjmN38aL6fFoTCJPDk7mB8URNBMYMjjqkEm8aYvo+vTk5RerBPXXm9Herww8dJ5uRYgORG7n+c
Nl76Lc2zK/TpQDLbX2s+gIpM8b4XkSY4LAW/zWde0iJPmM0C9aKXJCDv2QQx5N+0FZ3dUR4VAHJf
VjiO6bvHSLYDbzmaE9kCEpfVFy+jy36j6AggUHXyPT37ME2Vuzax87HrdoW1DV6YOqRjZsohNefR
itS1n633LvzbqmEPseAq14RGtaGAmcnSzKDyXWEQ2Nt4r6IEueNrdp1Y7j5xi1jh6a9KTg78Q9Ig
8XuCGiweC1SgK9FohxwAb7oLCbI0zvXBUKB/KIyYj1czx2vI8i2Hsxb7I+ZXE2oZi8bngvARivmX
uOVHgRBv4StsaIN1/9h6B6SANHAd++HHKXWXegWBaGw/abVOlcSORtpPKvwUace8z5QKt+YWwajK
W3KDniGBboWzBCFYYBXzxGW52oX35ZG1hO1pBMzvPIls3di7jRcV9+Q31k2SazudLsGeG60AXHuP
cRqZA+b0BJdGVxZb4+RVfSTQD7g6BhJ89+or3wfr1aN2ikpWkUAbY4J+OehHeFVZBJiMkvgdvjY6
DlfNr7L43Z7tgORPk3Nf9TBvHrrgAS3WjoFoP0LcYPqKQnl9TG0HXDL2d8E5kTBIgItN2G+r7Ke3
G09B+crmW1HA6HGFhPZXl90GCNYYah0EefUT44MRn6+ia/3JvfDL8HRq9ok2aZwwx96wAJZvD1aL
0On1dcEY4U9x2nNwMKcS8GlO7JoAD3YGPm3FHYV3NCtA9KgYoHLwNZSgFaKq/6VnRtI2mbKrZcKJ
E9r1cg0VhREhfrDIVNCZTRNF4l9kxep/JEO2UaX/MPXak2kaf5Vb8eEe54rW19NWeCkL6sx9ojgC
oVXgTtDqmnnWqTVilqVunaDGFrYAP/o2WuC97q57kgsVJ80NFg1coEHGrUzzEMsTZLhcw4RZwlGa
x3gaM8RZfUR5GjCc2pc33JCig7xTAF8vtIa1VbQqHIKqb+ErNge0q9vjt+hV7aJKCH/w+Loi5aB0
l2uZKySStVFeQY77/CdKvNmhNZiPztjuxoB6tpCs8841os5kl2iFr56ptyBV3LunIsgCsMzlKTJn
pMWvXvaPnror2PiH8GnY7gnQ7hlmGtPrI+MwKm0pZmQoXcgUKcyihowtb5cbiagLnA7iY5kSs/gU
mnJj5qPpMwy8E4fqezXfaVWLzHSHMI/A0WjRpt1BylNIwDlC8L7Lah1zKkzilOtZksLit7gtb4pU
V7jiKePyJIIJJfo0ByonFNDoYO5Vd5SpHvs5wMJEYJFUPbiFX2kaqKcyZ8whT0/u95kdO2fC2uU4
c6KYuUucQpCyVBlfW/b285dKMuMMRH6NT4xLOj/5uiPdKq2xhmOvznct7rJMxLORfm66OkpXXxKi
L/lia3q9JLrGWcWRg+dDlKI5er0sLCkDpHCmKWyrvIu+MZ/okCn25mXPA0xJAciBCdJpsQUh0UWT
Ga9BykzwY/71XRVjtS5oDFnIUWQcxKLE/6TPk4wBWkElbBZufEfErN06eJyvq1jZZZ6kpVg3vydu
y+CT/rBaJ6ByyTt7vHBsW3ZmIxO/XLNI6BZyl5RVelRC/GY//Xf/5zb9cosxU7sT/+j7IRcn2+04
eEzeOE6l/NSiMQ1vI/SGccX1vU61aAqMfHR+JZfmWA7Ow9RFLoU8z0Ymh/E8v+dM0uO33Q28sPPi
rfrcJKJuMAIwWWN8vQyYJ/IQrsulBiwo9lMeB+svffYnT23ok828ms3pmmfGJ/QREetyOoTnb540
baLyLJiUwxj0HPRRIXrH/gcgyVfVmBvXsNtR6S/55WSnb4x3de9m46esJo9tMYMWOfd4Z5NTfr/q
YfYitiFiMC4t5Fk2FNwoktiQDWF3pbpAa92Ej8swV4NzfUXez/TYYVERk/MNeY1rpQHSNDWsZhFv
0fEi7a8DVvge3PM1SlKLKu5uG94cIrpyywgvQPyTDLWeCzWcq4bFqqBmkQRQl1WIC8E1GyN9JjEN
PZKUPZx2Q6VA8b6D1Q549B7caoDWslWakpi5kdxC+1pICR/5BCybxRkoghvtyDg1d0VYXNdzr+gr
Keyd5YhmQ30herotVlaFzeCuuoQ7eXIJwpopfgNlY+CfnRzyIgSsSsCAO97IWLiJ553ljOxSSKq7
I3gng1FFY2/daCG+PX+nEeoZMaXGMDvjZCSYxzBYaM1wHFIKWoiLY/j4Wh1TnztzjzRpABcrGCU+
RQ2PyLDOx+GUoMSACEbE+rO1p5Nbf2q0skXz6vFtiWr/uZf35hL9rdd9wdh9aXSNNJ4V+C90SJrJ
n/lpNOXbU8VjWpY4rwrJE4eQjSzEmakeMf2RaY+1hIKD24VBKJOQ1arOu8nqkr8h/gpcYIqJAJVX
Nn+crObiGl6qvQHWkPSZO63vUnA/RgBxkOKAFRrmkd0edxbfC98yFbBlguiKKbINiluTOMrPry15
c3q890oQhlwQDKxGdO32TeGpUXBDnFigDB2ri6+SodjQPMpSy4MkpPoA11CaN6uUn74zmdZ/bAwb
f/D2TGWB5M6Q25eqZk97S0L+XBS98r7PQZQWGTXb1KHruSX7qbTNrtxa/rEldfdiUd+E9Ryzzb/P
Os+ZNGQ7ke1VkZoM7mJHQ8fVXUOLc8kh/7P7bMDlPbxuwOZzkpguoYQ9g1GSXg6VXgkIq8Lqq3h8
/XQUoVio4dZiRdA05EE5lLLb2xHmEp2CJbqxa1V+ALdbW7vJ5Rr8O7XAhA1EgDN2MWyPfNskiCY2
3IhRSF48SctwzqcGqmEqLoc1k6WzmFiFFhAOwiFy/KmKz1tWb3BOzF745hZjSMbJl7lJKUT95ZrP
ojw0c1o9hSMCwzjTp0ooj36Uh8DW7k51f4Pp5mmsava1noeUabpTXgj2nZ+IK9eTYj4qlxjM6hl8
DeXutY1Sj/4ZT/D6sitWIPiYVYOBC+o3KTroGNGUhCkJxQ8W9iNoZyLmCX7M5Ss7tv2WpcgjEjy5
LltvOIEBj+iUZ/9EmrOTy3NtnNPRg0YAs73Yvv8rRsRNWu6+MqOppr4M3PvpKSYkduIGH9AXE+H6
VeS1McaDgT5zkPndP6O0UTqR+HhGe1oEl4Dn2z2UlZmj0nNclaYkJYeUuiHy/yhbdo4kMVqUaYcO
tWvNtir/P3Rgn1UO5YXTkM/kIuuiiJ+iwWuq+tDzDlfbie26xzDgxT4DltZ+RiuC1yv8zuCgHIM0
mIUV7GyX3ALHq6yWfCkBPwFPv8Gn+xLbCPFfN9xh6075+uP/ZS/XSOnuH5BgWvbSW2ukAxFfkrht
IvZULm3tHku6Rox8ioVO0AKI+KJoU6VrRhDyKEJHh0B8Nlme1BgfKf6UgtTaBMxLSOjjdS6cPh++
ztrn0FOWDfqoPTnmrX2DEzQbc0eQo0XmKf0CTudyVeh4NZbbSYxRCQEwLAYk55Yh0bIQO9uC4hEj
PIVFN+C533Ga1AHKsIpnpc90iPKDUEk9tGyf0qmkEIh4W1AhwksWxDsVnbV4SDfc3+VOhl8SAr8y
ZA/oVPORxisY0phLhhlLq761Hw2goCwq1aGed4gEuKv/d9LYFYoYh58S5vuQQmJThgQQys+q3lqB
QtT+CIfzMzduhlmuN+O/5iLumFPZmy7RJZErzJPrc4oODMAoXv6Vo0rN2zFmnwT93Tw1HIM24tCE
n6JmPrAsDtd8i+yxfmO4+eNA/BZjz4qaAAIQo62e3IMFHA44Bo8t970fWH5rG42II/vSdcGLKRB2
H2PooEO90Ld+QHHC3c7wIVufgF6rDEWJIlHdneJcAOJoy1Euq/6T1qMvUwuLqBTiUT87RXe6aLlo
ZmZw83jDqLGNnjD3ImujiButtSBB3OF1tO5X745ee6TcF1Z+HudPtNLretlv+VxDNrZIOsInAVG1
I+pe4RAgu3EzZ6y9VzDugrBkiOZoHbmFaaJ6hhqtIEULnlhh7j9cC9HtR79nACEnPSG8q78z76HH
LyaeFjdYKe1vchDoOhoIkz1smyvlW75GGoneK6FVlOolqWCKO5UVfqX0BwO39Zo7ielVu9f0LdSL
rgKhpIFf+pCnS4gXecfLSZQBqGBvRlj1fwQwxkF8z+IBPK24LmeUM5DcYeuOoIU2fQEFIVI5Lz1z
knJZppBBjdRoa7bxFn/hIJScTLPOcuD0UGUe3L8trFuIFYiITk+zmc1q/JjPu66cxFqihbnTBs3M
X0rIOsP7fd6gWPGQnv0QbFHgaCE1vDKi3OXBVkiLng73538H16XM8ZLu/ugaJkO3Cgu+6U+BtNcL
5AP84t1V7FNTd4DeirDXHpGO4sW2nwFSwPhaY6Q+EAjvO+gAPShsbbFmUhAUyJG6v+YGGsWgcKI5
OZChPOga/78UYWUsyQjlAos0l3qWe9lBU8v7W5HqJ1DN8yWz3Bzjvot41S3MMZYcxo//WeSHy2P4
xzccxFIbJ9vRTUtzTWxMhqHGbc47ZJ6GRp7yH9o454nj72VFwWH3XZgKWFana09w3abYR1iW7dYJ
wQsGNoJsr++nMi5HGzG2dnNpN15YtYdAdIQQslYpzpz5fXsovm8wrSX5PAE35bxN2D47T3dUM9L4
64iKRayJX1ZtgGBtlZibbVnTrFPzg1j0xTpEhlWT+gqpDMifzLjoG0Cow+bQyA1Hl7YSV7KWwzBj
r7TmMhD2RrvVoB2eJY+USRAv4A6luhgGPC0wNxdz9z5ivDz4GTtC3pf7hnpKlowfzCOSxrNGolD2
N/dhRPfFpyTUJ25I+j4UrFnGW+hzmBO4Lq7UXnwffIZ5S/K8Rr+zLzPsJx4+mKdJ0BLztnuSNTqZ
avhOrGIb4lYJIrWZYM73FWvrn4jUEeQjIBdVGdTkz+2h5xwUpjtfKTnZsQmPoDvqdpRjTCt2X3JK
Inci1yydzh3aYMYst4MiEWGQzLOLDdMTguprRYiIEW3Ph7OW0mE5z68A48lC7IidqXEfvnLf8R8r
2cavy/ICNzyGqXPr/QvjWcouSDAPse4ZLNdynvBOZhcTZhoQWYRpVa346UotLh/uzr96w2nRpu2i
LsZt+EtCuuPB36V90YKQ2NL7xBMxRM4pVw6Su/qK63GbRYHK5vWCUIL+0nmfoAVlmLb1bu3ZeDFM
UCxgMfNOjAojBS4Er0/fHHlfKAttTcVvNFUSEDJvCy/Z8QuJ9CBCBUN8YUgOvsYhuZVQWnazxshd
P8d0VvAiJjymjun9VwN27vYAKEZzHUArRDR+4eiDdcRBL/k26JCJlmsvVEs0ih3Q3Bnx7U7nVsI6
g6NLrTTylQZT96u87e9o7SHsUnbya0u7/26Wg2InmCf1VKoqL+D+VR7FEwRwJdqTTIRsd7taWnMS
gppoAW3B+ZfBgpj36yP3mGK2D7JdY1Ie/G93ZI4DRaBOhJzePIQy7gyB4Bz3Hv+ToaLP5zbifdwx
sPsemnB2DTFJ1x1S+ly30z3aQrhMETWlSQDcu5VXqdf8FP2C9YVcjSx5XmuhvrsnfGam+hGgvK5S
yNOU8RICQ07qi684oZ7n432BJZC4udSzPmOZnmKPfgpQTVtfh/YjQVONGtCfhWjAb0vLdi0jwNXt
iv3p4NVFAZ+/OEqSNslBIqI4CSCULnXzkJBAn58zZVA1QDQrUWCSrafPgn3K+cp2aCx10/FjcFUS
GpsdzPVhyJBhYzVnoY99EX33W+NZyg5TwrLFscTG/Y44C78nYr+JdEsDzzg8yLrlKOmnChQTIR1x
xg+TeEHQaRxsbqovkcZ6xK3ilF7jI7/5KzFdAB+/jX9xpWs71qmxM67X6NExTh6auDIiZ+91xelw
p8hBg1RO9t8FCpdattiPMeCNry3SejIYANmxstlMU8ZDE4oDcrZ1INw30wTyNJ3HyAuBz9lTM9MZ
MdeohED4hNSL8ZS/98I6Di8MsZZV3rurqyO7soQNSw6dBk1FXdab03VPbkC+vXGvvjVXWw1k95yP
VJhibgd+6I666+VnqANoYyZughMb8zqXYfHv5bZpfM49LcXEA2RhMUHlNVKLWt82XmiI2FsMq3fy
7wetsMyw1JL70vTX+kueoaxHUQ6uxCWFLYDGY9/lq0gwtl4Zf/rLng48FFG9XGm9DwrMwBoCx60G
C8IOh/nFgJoDoLOXEOyW8hBzU+P5SnhZsUOBMQytYXNWYdS2caFyFviekKKT1OYwQs1ozd85CwCo
I9xeA6M6cV3eyych4IPYdiT5JzVd0AFKBaVOzjI0GPd/z6+hS1T8tSvm+j8ruHOGlXhOJl4/6XwN
GVFKFqlWWTxA9iDuVMOzsdo/F0lSo4Ur8kdJAhfVlqTgfNpWDu2c/V8Y66k4lL7w+49e/x2cNCsv
vE0gmsR5wOx7MGx/nioZ8YWI+S3wPFExKl10/+ujTGc5gVmUsamAd++yFRxmNW1t9QBs8OZj1Q6K
nB8Fj1Ar5KIOBMMBHVIh6Tg3KaeNEJ36O7TaghKnembZNDqzxQn2n6XRV3MHT7OM3mThRCoo9IB7
IjhEFOtFzZxmuVhGMb307k8kSkghFKtDc4Yy7kU9SrQw4XEike3yuAx8eGZuqM2tswTXPCv2aBiw
ohGfnTsfBknsLsYRhsRn/HBtM6ABguHXZb2Lc7h1uVadykHv0yQ+R1k6+uhKCiRaO0G5H2AwOUX7
ErPXqeV/lymVikVO1K72z05J8BaK4dpe5MPCXlMbjmRNviHE6c5+WF8szDIthYVQ3lDUu0DZaoKY
XcQvLX0pLftd0ggU4K1FGYcZOPP6Qp4BtpyqgsBPMhhOgOaWSylWbbLt02I7Nhq//AoAQqRAxmD/
6PzCee67Er1mZBLpzEmmTXTJPy6Fqxb10mftTnO/K+Y/5qSpbMiJSga+LOo6SaoFv7LDIiridIuo
iQAMuK8pwropAdxOqHYc1k7mRiC1hFuz7rp7OI1Fz8ZnvTw/o2pO04Fv809NIylYUEp3CS6filXq
IgOPvaWa6fCrLsnp3C2+UzE8kBhOZlMyoAcPeNvRKCZg/4n1p3m8B//MRupSNiiUX4egrRu+u0nb
qrxy7v378IU6+sfahJHLzmFZdQQfXhsRAPDurIwIDrVm955Rf8Gvx0V/k9yYdm5A+fSrSfq8su4b
vB/W1XCDM4lKjGmR6mWj5eNo/ae+FNnc8mGIAdfFRMm7EoVqn1F/Ms7uk2QQ7fYsM/H8duNdQH8g
qfGDBM6a+uuILaXHdLTk0WU9NfIf/e4FNkt8aWU4iEUMwrn5bPA1glFWTFpMkMAH5amK6o34EIx8
nGeWSfEgZp0FZu4nLCkOTBzQKWWc7MapDkqn9pSUiqOaPTvNWehnQWuwfAYQBrgOv0Y9sR+M1Gwx
9n8ZH2kcjGzDyFLR/EoPinvd9NS2fLXQZXDJUbOjrjzbe1QR7jWgBXhhPi4DzKA+tNJ6Kw6Krlvn
olgbcK6llBHWAv1YxifqamyJiOkcrwdHcd7N7uxE7KaBVkt7SNlHh/OQslQ/UdlDQ6t6wqnsI2xh
mvGXRk2hYLBu32htk3YuygJPxPdfsPVWgAVYA8prV1hKZt58EF7l+eX7Sbfuor1QHRcFIx7ljsDo
IArzNNiuq3Ri3+nml3RrCif5oce6bYcuwFdI7glH1SLGLytGJCnP4aIQIzGsY0SO+T9cc64acgGS
yysnvm7SZ8X3YoTTujUHf2NQFJWy/89BUwPiojnbGAY3CH/FDoWUNhch2exTb/+9fuYSzKbpcSA8
sY1IB13a8fKGaun5YG+7JPnxmx356IgIcYHwE5M6Mjj85Tfr1i7v2AxhxNrFdRPPR3lLWLRsFPeo
5fDSgEdmEvriDiQdOFsfJ0ydA+dv7KFnp63bf3RIU0taPhOiMgkCAAz+cWVB+tTkSqPBpf1vLO0U
OoLgC5AC8w1krz31TplN5JP+VsHo/4SbZRdnC1LMgw72KmXsVbwsUwywgpaQtcyCIVpq3CACtP30
NNegwdjxAD2PajYE3e8YS4s2dBJZCcIoUPmw2pVNysfLow9SQ3+LC5UCGfzOUrnwla8nUBIVN0gb
S77FysCYPa38C3tIKsM+/G8J2qE7vJvA5+ucJmOf4bZ+XpLPRoDPxCSkEfn8z0JVcaa+uRvGY3/y
JF9lyw2hjtmwSGE0YRTbOOr4TGCEkZC5QZRAYH7OxgvvRaGxEI9pufRg6z3LdxmfNlgXXR0NBIIa
Qv0La45hwW/J7gwl/Yv8fhOAbjLkowin50TLwWGI32Oc39OwCR5xJ2OPZX3RAuVsENfZ8PHxyyZS
6AlQh1drq7fx+39EuC+MxDIPSpSeYpFljdcLdVQD1zb703BW2PEeI5QxIRZfFi00wBwQWuwL76EC
ag9YZleGrVrow9wAkhdbtDWtcstU7O2qUVEa6ZQ0DJz36t7zK499pIv/mSxbaaDCOakyjDaAeJzn
1Kgr+0c6UyDDFyuq+9dytE5H+Id1en7b8ML1/0qUf0mzSZxNW9vivaMeyUB6hqTdO1mGXIFjp7n4
7Ok3HvQkqbXoChA4iWSRQdYN9wwUdiucpTPDjyhRXIG47naUzUyKLCVraVA3vd7FEwteitDmQMgy
39/ptkX8s5RFn5Xe4RrQE2nVa5n2I+85FAL6NfHXubXe+oLFq+8Ef3p2Pd3iZwm6n6AGe3FXclKt
gInXwSkFMgs1HdAF/4r/1c0ryktcMpCEVohrhRh4y5nbH+wCZwqYRBxkaHpqGy2R4z34HrFlCodi
NEP7NXo4qMWAck24Vcm8mMhVFOrojAYyWUACzPMwLVBIjEzK+3HEOpwyt7TcJuwPv73G++lxte/k
iHEFur3uwlDQ5FGdIi0G1VfE2aGmH1uc77EgkYXdLk8bCXMd9O/egFrLXoiEnMwxcLnI4kCsFtc8
vh4ujSJ2WYy8O8rg3OOZ6esXP2p4c3Yvl27vZMqv1yIj4HGEgog6OLMLX8U2x4I8TVZQgBSrdScr
SF571httmIYay8661NShv67GW/9O+y9XWm41xqmuvVfooHv8LMgRPOXOF5b9bn1om5jmRTiyVi1I
MbhBSE4MSmZq6DNlli/tXMhjWVnmscNYAo4QWmgV96yxuJRiHl8u1oqZyCQvB9E8Cwm+AAViK0AI
3Mvflphnp4XLnTwJaVMDQKuE2LD/5de97LG5ulohsVkt+qoj57JD35zjnicNuQaYWPSxSXSx1uUr
ShcKehXwPgVTVtjm1+Ms75MOwmTF7L3Al7YNMFKYRF8RQREyPz13lPKz4d6ZP7f7LTPp6teItzC/
ba+0UlyQEQosiFBVzIdRgP6HdNiNDl1b8AYFqUybKNokhiTPlfjBpwHY4UpojGyCLPqzaDd+TnCU
VgW3eOlFUyH+HL8j/+roC2C9XpI8lMziEL/2V+uDzmKaQUqrNGoD+kXkY5IO154dDHMMKarE0QPl
dY2/wVCb57oIzyaPEP6YvVoeZzBstFfPzIdGKmlLZ4Id/b4pzchs64aKYfXA8b3+JFswzfni8rdS
K44tHK7Yf5svZE9hy4hKu0FJEzI9H0X8oNH0DTCCrIaiB/ifa5GLniW8idMtr+5ehcoeW7ygblpC
SfwtSxUI57xY21ALNx47r6W4dAU04pWOsBg0WTImGdn2uVZx4Udw3qLnwnfnXKSysPFNlXbwuAnI
pC28kvrTkwJX95nm0VJf5FpZD5YTosiJn1gKgTAfSKNJSsPyzX2xvBhMeRvbYrKKPhpKqB1iZ73B
ZS3ATELbnGc+LMA17WeHytQhstA78X4rR/etFCaIq0GvA4vJYl298M2eulA8Qfj1s+oDD4T1INd1
wdAqZp3nXip9iF4ywKVhze82VRzlQ7ed8tJ2XwpE5d++KsZae1idFk7WBQNUUc5E4nZhB8JCWO7m
FPHnPRp2McUDQIkckbU7CcGtPFN2zY9XJgciHAwg6O6dZa1sB2Ef8uCOUDs3xiSsnZ+OR8Bk264i
ZY7SQykTdUcoFxNw+wH+oVkpry56jXKAR/XGIHSNUbe7EayC8sp/zScgdD9HqwdQQqdTANqXwQKb
SjPTF16z9EEIyQGwh75KtK5gigJ+1/fCx5YfDwXiqZDUGz8XEq8jlayOT4dsR7d8WjDrI6WXLGUI
LvLmXeDScEYOphnDvhLNxEiQaYa9OOl4jCGDNADWj+6aZx/geHCeDbqrv/UfvxQlR9VEzx1Zl9Vo
FEMeK4XsRJYy7JfpErj/tayCaokqWEJlPgL7jde6EbqdMcFU3+3u5C6/rJqwtwPHWkfB0xqoFenm
BexjasZyrFv1Du3NOnhs70nVyWmM1HVdIhq5sbw05UWFDhHUR46TROWTiTJ5QEYkHVI05P/y/QSx
mS8SXKDtt79aNtgXObvVUYbDI26W39IjLItRn4C6fiCFcNHMamtqmf85YIhxnOoVlSkH7LU/bMgF
NfkqCz4CH56oM71wZ0JMZzAiGBgc2di/40FUwg29N++IFLc8QPPWs1/424iT3o9DMqEJXOD4qYgo
UpYJeXzg19NlYQ/ITlT7MxqRPAsH73CRbmU2KsLXP17dd4UHTSk9Awzkqb1gPQvP1VlOy8KAECJG
VgbQb7rsSLvcnfZyJlLQBgF4ZAN5Q9AWh94jvLO9K4Fm9iFSQRVnDu/yaLSMNG4MHtocwXBAbob7
Gpj38eouNFzvSv5bm7IBooBTB+BI178D2WbAB13PHPyqxSYZMB0qs0BJbZisJarwFq18OGkjUmPD
yWdfD6npNdd7DsgiqOEukLkTifSJPxv/b1EBGNzPfKwRlIkVTR0MRu+ptqymeQfJsRhRDqg26CNo
99QjJBVdYAJDGKnu03jSjnI9Kr2pitr+S5aLo8qP2W+jvriTO7eVqSeT3+Qmfeug9UpqF2KKbZ5h
e4ng+2tL4mpnBlDAZpeKbOz667FGMBDsDQ5d7ysHH6+m5D7r2VD84RJw+dcg8EUBZ+1F2rERGE9f
1RzYxH1szzlUnALPEotnWenRWjpTEXa6KR2b0rofZ/9YCfqnRUlk+Idf8UdGZlPwRZQ3N8SagKbX
N1w88kMvoyZCICdn9awJ8BH1E8j2MHoUGXNP7/9aEGBE+ISWM57AnZrsFgzSc7NtNtFjQTtSLZv2
NnVSfFHw6lR5gKwNVA8giNoKspe3rfXAlYn5WRWgLEmhbVCg6lLjHglMkX+OS/annT/l/wCt8Lft
UQNww45VQ3i7Nixtq7+rbC0vgEB151rf0jZp77PfpEm9fI0FXW5M+L+hvuSkFkXVN7nt72SsmauB
Ct01b8mPjc9a26R2HWcZrMcIL5tZPWQSY54DvgaW3yp1qkh0fAW5dNF11MEqg2qoGcyzcp7Zpse4
koTF5lyVUG71+iQDizQHXAKLIoYnmbPAmkJ64EFR7h44PEqTqqxTbcgMHdVkiaMYhNb+D8+yUPeH
MvmrdOtJrx7wA9jKfVtYbd7/Is+wG9+tjBZ9fZeGCAwTKYq+gNR/X2lqkJcxCItU62Hyuh7iOQyc
9McCmZmZRWA5tKi1VeOtDL/NXHNt19UR6kPVmTUXh4IOXJmKOnMQeW5sIo6gGSw6XUN7b5771Kwk
8UBtwRJWut8H37FaSgg61+fIMq4Kzwyvb6SUsXkNwRMeQlZv4JbWIKeVMlisyllK7itn3rImA/Cg
3HceEZAR1Xfc1jjYYv8wWdwgtmmHA4KaPVWpo922T+6JHFvYYEv/N7lO2IMOEr0nWRkdGb/jgPaN
adfXNcahbbNDr4oHHrTRRq0aFK1XEiayfYxOYNWjCQ4I1CrFNTEWSjpAsdXZo6tFVPUrM/j/xuyt
hN4Ni2h9diOiCL19hElXqacPuecNIuMBXS8wkMb9s1A5kSF29jM6htqJjl0PRad2+7hdfkRYqiFm
epYhzprUAQF0gg5G1tYTgMXIPJQQA+XzTG26THdjHLVXA9o+FEzMgI3Jbdd5ZR8p84vpkT5Zba1n
Pw4EQm49RXoWhIXFY9TnJWGXsjXluB0VF9lmnQ39S4wnARUIvdHp2rjOJzHiGDHrEii9NMTJt/S+
1rV1bmpgHHQRz3HSqbeisWfasIr5+evqq2Y6MXq2dp/qHnjJdAJ6MqS0JExtdoxiz7n2i0SdtVSy
sBzspGGGD8OykNO0s7ViMlXJBsD4XXgABbpTm9TcoGnki38kCJSm6N9BL30nV7PFHt765NBvA+P6
SGJAD7uUMqEOUxyUlcxoE/tioWl9RkHXMc8FV56rKQY8JMSDR8YKjKd/B6Ap3/JZ8ClBdJyDqmzt
umfHYEmCWobbbk/ZVNUkkLkatsO3BbGYKM4Dweto3bfqdntxpwkqi+v6pAB76mOKdO2oupsy8q3O
KnqJBuC4dd4rk1qUUPHiy0vY+9PkACRsQ42yad245f+lqezb105Nl4iiG0+NWxZh9CXZmvNVlL5O
dVBXehgAHQ5VeZyJYPRmxQcUT7dsUpzZY6au/z/UmnQzwEoN/3g5+r0f0NZiFUPVY0VwjllqlwUK
wTHy/PdEJWNT+A5J7cMtOTGLps9Md4iQU1oNoKF3+PXGlMgGgMid2fQh9K2zC1tduGxp09Fe8XRO
QiU5mn3NQCJgUtfP3FG7dHc5G/xwF9QNSuwW+h4ZWA95jjDGRfC5wsgma5WNUtnH3346/24bouE5
x+JTZfhHuDmWc7SsNNdRWff3mN7U8k+9Q/3US3FzGmJXgz2wz+mFrA/QhSOQ7N2QEwyIdQ0Sqy6l
sfIPeIvSx+rEuYBlyJjZDv2hwe12VNdmfoT6NT7otYyZXvizS9UQfEdC5yL04jj3T7a4YevH5h91
q3lWpr9nTG3L5n33oaQEvcfrdpU1M+1jJU53bQDbEkXX5jhJTdTu+xADJI3AMbZEhHDNYzuroIR6
o6eXYw8zL264ZSq+ZBZrQAX2tEfyLvUw6ykIWKq0pomb5j9aL8oArgx3zugpCitWCqx7zt2fjmul
woOdtNJKiIv2OPuHHwK6vQNu8cwPof1qEOKUGaxaB6vHX7LI3JJ4EL0kwx5GAyhsc6+npUC7/jGG
ouU3nXid5H84oJ4Ae/I8Pm/o4hnM0BCMYDZk7P8WYMGqCj8fPfPuyGGG4dishmL19uRh00JngfYL
cbCMj2TrpoIahVOolx6uGqygRNWfJXJjGIwLWlEgXHGBB9gleIKyjxnvp7ixR8H9z28qt4/TMSah
zBHeFS2B0B3v81/cyZnA2Kf1T776I46e8vhJVhfC1o0oYh0DcUS4bOycGPCR2TkFK/v9wtMINi1B
7GEybzcZfQE6uF35YJp2ekM6UZxH8VU9CUqcqyYjrwo29OlUc+78YGxu9vEPNRy4kjPLZoUUWfTa
R3CsB0T6ABjKOxMhnwO+VxtinnawN/zhx/c6tvYbekBXUSi6Ei3tf5YxV1qT2lgG3VtXVCmqwlK8
TyoYWLnJlqOqt7qrBitdmSI19sWBWv8Lh/t1HbqEue9KMHMGqJ01/9DgqJxrJIt4avVWK6vM5jQ/
paoZZHnun0DjIxON99cQSt43IlbNtssqiI5eXCyUa4WHHmL1BQ85z7co1S7W9pXTKhFqXjR8/Qi5
a+lCCNvMw7fisNL2hsfWJECB3LcNvZO/Y4UlhIaq2Zd83EwjnyYWu5XETx23fTLiGcArTaoyGnI2
XJUsBm14J/cWUZgwUab2nhwk12DYGaYCxCJcDDJAizmxmxgFOHMrp6nWee8a/62xl84790QzB/b2
IZ0QTdZP9E66nSwYN4Z7qn+/Z3elrJ0JMoeBI4kuvhrermU7ICHIemRaPA68rn2+ovrujKjGwbh9
vrBWPLd4Jeo5JQnL3eXuOIxWY2/OIjmZ5xs7CiKkAvGi+mTXcTiB0UEblxh9SkIfwbZcvl0mZsAx
BHNhqj5moVjmTZOJ2Wo1tC+uXlB+GvDpLqXBq5ZeUJFTWWNzMCTBQtPj+9J+4hjBYIeaMgXxoOWv
vAzTx5qqpBeq/caox0iCopNvJY0fvsvWy7hbxFnY8aaSb9H4knhXhy2/KRHV4NDy7AsVlspbiwdC
x566Svesk4WscwJvH1TPNIqOtvuohxaXv5Wh1Nt3I1hH4ktP8ZmHtjeCMxRjOgnsdiOihf85FcPO
s1p0H7/eKk7VhcVsN6v/uwiXVbQFxjiUQky7TAO2543w90SQQCH5AL6LpmCElMGY3RUMyqD9kITV
2PddQB1/Tpx/uQRxZFdCAHXQEWHPCanakRE2G7X1q7zcXuoUylLfmkk782alufW6pkw/iDVvlpeL
NUiqtzsGbxejOn3Gi0x26JrFuyWzES38GTDABI2OczjqiO3LRCwZXYvU14TZMJpm9ZMgbiVJLmFE
oDSo7Edz+AOQAUpuUgxyEXD1UCee+ffbPe63F5gsHVsPbhRreUF4A2h2trjJT9nkFOJ6IF9F3Vkx
DwS5D41jaw66rbfRLrGi/GWmzBXdH+IfMyqsvBmJR8HkPwRGmjnjOAyj42HHjJuQ/cBGNkptdC7H
zwl5w1mAOWLmrbQPruwcVJL1Bu1U0aQ1CgLdp8wCAKOsnmr6tQC3fY9wh67XpV+CMsnVXfxQgqNG
2/Z9aG+5wrrbU4C2m3ZzwFxeIGXvUynwpNU64rgDb83u2OQx9CgIc+7v0iT9SvN6voAlzShfDLxE
vGBqn5qclO+hVbQfA8EjrOooXCcLWwIGC4clILJWjQ65wnWUtc+aVC3m+uv4ot6AmI9a1GyZAKUM
jaOMrWna7lCPGGLnrsTZBzx4qKgnFGvCe+UeMF1GO8TVOqCNa9QgVuDyFR/Q4lnrimJ4z43kz4yF
zPruJm4LTncePVtGY7zePArw5AJjhrN65O4SRUQzdenmWXsHAWLNhYdmjlX7u5HGIkI6XBRn95jU
/BG4UXpzblSqjpxXShIC9UmrPEvWtUwibqd9+e4I9BYPH+8+ruYjhjkT3P5r7z4662LUJ/cmDC8p
a9UOZCFcWRoRbgjWQm4o9QtkKbZ0cfaQTQIxjOgdJ/kOFfjuZdcQW1/j/4K9zXA7nYkwgN5zKgVr
21X1GnfG4xwVCRWY7QBsy8Oy3tuWYhhOFd6zHpLQhBRsZMEjGHFJy+YJMBhb1GWQN1CVqVsWTFou
4Vhgl2Kyq2RlR1Cjn4sD3VhsIQKP5ew/0o6vMzABYCGDzsomUaIocAy9ussGXJntpKaYo05Ay3Ju
cyfaN+QgxfoYBCgUgChdX3QJebT1ZOcscYbMJXpgVx1uUuZerZIGFHDtufpyYeEnqTg8V7PpZ5Zg
fqVwfSFB7AHGgmyJXqjDiMS/loff/jP1Ye/PEZfB4xs99aIYK2Rwk1+i2r0TtGRxjc8+YlNKfn/o
Tc/35nQGdDOunK0xdWEoaxLbiu2MuTEeJtMRMW6vS33VA3cgFh+zcLj6kFLXumnsrSDZuKAj5nJV
UfBqknpLWSJKF4ii0HM9nvxdhGpkNYR6zMLRUrsZfVkoyfD9IOikxPKT0m4PdYfDqvIbVNBsO3ql
0fmgMyWP8wuS1FdTSpN0izl2n3+YLxLuESpineDc89CVuIZ7dHhl9oi3Hb7UaAGoYvnTnUP4xTau
GRPWZ5pN+IqQpp9zuSZGmwtDJFq5CTVfbBDjCjrvZrKxz50s/YQTt7ArUyWazpTd/6tcJlInJ8hR
sA1PiAXSeZ1pJGZfmHqBxFY0b3X9v0CAo4n2cXOm8UnRkIFq49gai21/DDqmnyTQpAbxdtqoczdz
JYPNSiLsYoS3wh+AQZz2FvwCFCnywCxAkHJyFbcdQQZGbAA44GL38xrFLJUrRVCDN+EaxUy4xz4r
ZltGnNI6fqEejRCJm6P66qNuzTSyk31l3umi+Pj3R2zjfhDdiSqdNapUD5Ayq644crWHBy/1N5mr
uNy0TRIfL+bRK8ncZYZlTic8QeXP44oqICrA4rrqnT6FkIK5uEqWHK0FyB62mxTC6gHDirBT87o1
BXGAMZQ1cZkcLdcXXNBKVKghKvBztUtI52tjUX/2pomSdi/7dOjLiuC/JfQjsWoJo1r2e9wTm1Vb
inJmqOd10+PnXYpGJY6OaN/W3vUp9oIAxi6eEAcj8RTFp3ex/GP8fA9jrdoIaYZoThFXhYLM1HIT
JY8Tt3zqQrhf70cZjXXK6LLfO3pWTmdw1ZYBqVtI+dHu1x/Ax8NslK+MQXOej3z5Tl2TN+3upqcl
mBejqj3uqf+sthX1eligXGsZqSFJgWwwxjpSjVHqfkAYsvk2w3WgGl449/KrLFwZo1YUBcTXFLy7
ww0Fs/tf/ItZuOZJH14gq9K4n+fMXpgx4YNM+sxRmjplcqo5uxr6odhtIUP8BEsGJnuYoxiYHcty
qDh+dvydF+qNzmE15ERt7J6Cqj6PGLO6kCcbYwrCjEhSrYXysZKfE5sE88Ulqm3ZsILA4FCJRtMR
VrFh5qbr8/KWZAuBGdmlQ5Q1tVLlHqNypicJvVUdAEmU1H8/WQ3ZmRH9TPmesT1ciGhtkZoqtZO9
vofwC+ZsvW4LMFyboXzjO35AQjyYDaE3mHpJQvmTrPHy7DPxsVzMflxHedtWNXU13xsO6pTe8z/R
OdyBXFKOwDeSagbzqTx94x9Y39OmwPMWzV4g5D81aPmtjbZ4xQFYFGtvfpMQeedv92uJsnqQAN0L
GZJ2VO0tcHVJfFMzAmgjsSIr2Dp0y4l2TLQXP6cPujwz+f9qf8Fotr+NHzSuOBxkQNE816cqFo7k
U215lsLdF8RyQTwlSLnvMljTXxbLhvL3wQhSkHULXNmdREKv4Ix4irK3swtojfShU6Wnu78H5gAw
YptGwR3iAn9JRY/LF5Td6G7ylWCqQSPpETNN2zfjy28jPOFtky5N3tsy3iAXo9c2+ytGg6FwXfg2
z2ifwT9VX157MVqh3ejS/SDPxtWPaJE0GnBfg9iqqMSXTF/pXoP+XRT+H0aVI60TdDHLuq32QioB
GBaQnogcU6H8/KitYcuDOiV2dzsWBXRrUXVTeQyTxinsjQknbwChksSvcMg9UDeVylrThQHT5oF0
k9nCKFiPeeYesOSKvo/reW6TJV/duaZhPynvNphCPRAvoCTYZwrcWG/iBgrD5NiNp99oi6VLdW0y
yBaaYWy7cGT0TkrNApj4vK6yPq/lwI9ndmjLQdAuE5zKr5gbRYMevdx9j4VrFxI0b96WWowkRKL4
g272o+dSwYt03bjoW8NfhIEnI1mqtrTU0ETZLE84Wa+NebavjYA8iCvA7G3Q2wEUUVa+eEw1p+3k
Rg8P81XM2k6r0JtEFTJ4odwPjoDG3Lex1P3p8vsDkWoL4808bwpEcYyGL9r2dNl8hmGP877rdgaW
Nwe02uEu2OcCbNwgre2q+HbDxUL9BJzBRsCmAOzlDl1gP7eFZ37eR4bEtupbC4mlnOvi/RvEI3MJ
JHzWdRudgZA7Xaq22TResfHam1JLX+lkh+sr+CwBW70fc82GVlWlMPJyY86/ff//JmoBAsUMzDJQ
FNeLTMg2E1b6yeIyLi78fmJf2oZFTny8upns7hEjbBxQQ4Mk8rPurGAEqotYlcSCAkyNOfjab1zw
pQknjLI1/Wh12QjSMZa5mxquRVEezx/lCdug3gm1rIO6sY53QPrkSkaiQIqg0qdbCIhx6DtCl/KD
6vSMcl+GBVC5yGqwTdMGQfbTtf0wm8GAqSGnNc8/YW3IuwtNCmmOmRoy+UIYKVLM1drIqDxBF4FR
vwl5ZN74m6SA0JrkaqhcsCDFN7jW8mdyvhlpCSHh5bcFbL2ro27snA2SYvbKaBCIUpjjK3jfnUgc
TmBseix/I3ek/lBuR6GhLbwJQi/u7H8AxYBjgiZtlREnTcPbBewqYxm8JdmyzyXpC7FOwueCUMKH
U5lg7hNaU2iPGOQp5+zwDAYc67Z87xlBdxBriPzN+mhSSRQ5UqWmLBJtr+gVFHCEFkZgzqO1TnCC
UWbnIKQkIxTUSeOMHJnKjHlVJhWcBBVhowBKSRRGnfBbrKhP84ukKKI4vtdockgNOS6TZmekWkju
vusYV7GTXArSQ06rEUl+pc9+ZkYeR8gjA7bUdBdF/k+fXonqtt3eCFVSnKM73efyIk/YYiHwh2gB
KBTuaHTCaZWnmSYbqhoYPa96D/tVSfSQ5+cZWC3jr8xfVKjbOp7oRI6nXRIS09PuJFEo0Mym0jum
eSMtx+xcY2f42chr8Mq5pErAdKdbrxgv3Z+JmR5fdwmyDwFb8zRxNPO2rG8aWPMNOs5dr2BZkSGa
aHn82USruNBIVo1Lzk7hiUEDOCFawdl9g51RWgxkst8unHQqQpcTvArTfs6sgjcNCoQqoLUqk6dM
LDQ5y1uLaQySNxGQ9OwDjNnknT18dUd4rD5M0usfnK9uQY/6B7fvhcaDsEf4ZnzdEwFsEnzEl/ju
GHaDOf1YJsC9sDbD0Q57c6zNH7Y/xu3SqqpRloOMQbk0eDlZ0129KTIFfiC52t14vCKBzqP+W9BG
sBWBkDeI/w8Zavjx9smk2+KBOX3A4f7UbYSAAc9uyR/gVBa3tHT39nR7pRqEHEBnZnOOaayhh9Ra
m7wIdzfJQpI/3NkHP2gUiBNw/uluvk8oVsUVcItYmGh9RElTRXzxjGR4sDyo1eLRCIN0sdi42sTO
4G1KXCamkXQLUfFPibcWlNfNk7RXb/EqKE07tzOyjAgwitafwPJimXHsydrbhSQ3h6yyx/qHBV6u
6S+xR8Eb5W1W3bsr4hfJIkTwPcdCmFG5TTm33cNqqm5Ntq1wEDWP1gV2cS+Uh6Un++0IaVbetcVb
+N/ntYBpOOBPzc62hVfsq+mtMjF9oV5sJiIekBGjlqhx2rHsOUh/NJJi+nwQWIegulKzDDTPlAa9
5eh7EXbwfF+vHXNDj6TmlyxWXsNUxR197cfxJpcn+8Ga9pgmC3yT+FTcWbWUccCaXaD/0z5zRYXG
Mu1p0nBk1BuGBR9VB92sRGHaqt2odjH+diiFH/mag3Mrzw+ywSPoFoG/s0h5cd+UX81kSlfuKNh4
kZnX1dU7WZ6yTBliGOBcstb+qJgD43l3ng4JMC3er3rq0caOjCaIo8LnDKnj/iABESFHd9++x92J
IzMt4hvFRhR13tEwE5TvyFgPCIeqV3iM/SbrcQb+31R97C2eFe2HRHo0ROjiXxLf4TmH+PcNhqto
dn3SHTN3KRD7KjyhD1tENbMxYuHpsX9akr2CViIEnb3bK8SS8+oET7047GdIsbs//Yld52Iag3j+
Er+iAu6UO8u89kv3t/ACAqXaNYcpJ6Rwyrj5HU57oULufc2W9wRJ2w5NqOePZbgzBkNq9xpuWM3d
drvZBDwv+FUKVK0G5B1YAzwm/k1alNoHNvjvBb0cnHpiiO93VcD7YDuy0wGbzVxGf/Vqb+z0AJEN
bxTUyCLrbAEPCd8azL+h+XlKjIYBLJfM/msziD/0Tm+un6VUtpPzpN8Huls14CZrItXQ3Jleci50
WtVBneBqHQJmDtbtMlAY99yl9G1bC2ooYAiB/6wIeLTBe07bt+Dq9xdeuDdGZSQcQC4cT9U4lO9D
cy7/+a+c6a5QGjVV0hF7gVNruFPYaWvKAdZIWJP7B7PJff27ssyu5mdeNBFC3fhNOKm4SHaYEIDW
Ru2ZiNhpZQKUa5jiCXZ+93Ke9kOd13dpKA453w+WKJgdkYSr2b8LQusdfRzYtG2NOzwwfTO8vQJ2
A4QtkIn4DhQdCcGR1nRqzB0vuJxPP768AWWIDHwxAvQjrWqX/80vSAsKaRLGrHhNkXo+1jpE/tdu
lxzCXuAcc40XLoYVTJ66XC6dC+nsOwbTfRjlxsumkw0ql+iV48S2vUhAZPSiZWznOZdXF88mdbSP
0QmquhkdebFn8bMyDqu0vF3ygBSTkklzUUYPE2b1v8Fyb7+x7Pp8ZN8veXS9RMjPnCxq4KWO1ERx
y9Uck8AHUprJNH/aLE8iTJEIfSy/xejwNHPevRz+MWUAqMmm7UZwnWOAfwvMjCCS/lazcOOni3Yo
SGQOgZorMsoJkhifXpiLZm7hBu+z+BugPUL8TecXncGvhNeo23pVih+ZOphS8un+bbHKeGdJM9Kz
9JCPoLeP3mXUeLKuuWPki6UkEYAWKP0OFoOxXYHCWYeqOldyBgLbxAXIvmdrC6DwjD+Lo41hQnm2
CgSUvPH6SD6zFEsOeqWaBlXcdiAVATdPiEQNUpN/ejAwm6I0JexbLXQcUUBJ52DyAlU2+xoVTf6D
j+bPMbYtmy3H5sRHUQEgGgo6FHHAvXVWChI064sbg2/VzDyGJ5ofLzVFCHPPbVM0MAGnFvyf5sb3
OVLt2RGoXQXMSATtXBpjeDZlmmYHi0mqHMqr9lRAMjlZPhIUoSQ2vp6cuWDQ5+1UCQpR4RAuSoVs
ZABiVWKJ0TEBItriJ3vrmLI6bAHJLGy6hQjK984SsUM3t9naFnIsWXxTNwEirmvC1dEpIKgrhYdt
y5OcGxWaxPtuFxqlx0nxUxu1MCr3KIvD8kq6pfwneqhmG9xwmTDkiIvpGI4fWSx6pixSOzhPqHsD
xOa8Tn5qb1ZBIP0zEP7Fq47RqZE3InmkCpZ2G3xaIob6gOIWs3UZ94oknZlcbEJiSKcCk1cxUmdc
CaMvvQxusBErbmxn+9jvTo1h7+JF8LptTrv6keTExZmfrqHqayOQc/ShehTmbfE0q+tYLptrdERf
pQYTcnx9+FUp7QxKn4euPmnLsQGKwglDnAfXgimAveefacjT7EzRkDP2/AFVh0ZM+AZvHvJnXrPq
0GDkptKU/Q80Plbfve6PZ0ndIwtkiiqdF36sZORzFMqaC5gvVI+/u8FH3swhordXmCaL+9y7Ig5O
wj95QekryZNDzJ7KRG7M8DPNMEPaF0BS+UKt+j45jsgZsQskJK9s8dRvGud0ckAUdtNnvSXGQmlC
2tX4BrJ9KjheA+7tepeRDERrW/WiqXhPXmv7XhMjgCOXPrfy/IQHuTkaJNB5J3F68ZRDqqxqsZ54
Ubt9uepxh2mW/c7OCWKaxWMtDmpNxKCdDw6zgKPSFF+ot8nSCYEBflyiNRQdVPba8DPAF2qWqTAH
KUMc2pouZKw2WPa1XIMA7rhjX69eKFETJrrfFuuRDAC3hq/BHyL6ksfEkxx/DKY+kZiZWQz8nASf
UzB/IbIscISv9oma2IheFWidQM8OE9DwsP8MjvbStmrIMJfZPDbdWvNz8SpUZvqk5aNooiko82OZ
d/HGbqW9ejtgsoQq+3xNMrfrwfG9eoGJxRe2tjn1tJ9Nkcv4Y7zeztGd9JS7EjGxA4zVP+VHWd0N
A8TQMHmWvcPAQ3AHoM6k6EdXtNFVubySjfmzI3XcaLhfO3oVo/W5aJ4mV9y3PSgPAeun/mWvlUa2
UfV3jgZl7RL9uVzj8mRdCh3EsAJ5GjiAlCqBa2fUynVsaoCCStPTbVNwcSFNX24H0mHv/1cVd3KM
EQ2qeqyCJWffEhplSI8+RnEWPc2wR4Tbzitt+2caZfNJf7voVAkpVvVBiMnGTxRC1huAQ/PA6JlW
Et9OAuX4uPJsa4Ifk+R+rJPdAOlbpsPYaqUAFGY2SgwEaiQFSvk3fTinm2AGaCalPDljigkeDNtc
s4DDI3QZR/zDLz2Gm+e/Kgwq0nT6mF47EYbmb/vIG+sQ2xsf3NAvCjdsIN90oTUESsMGNWgPODFk
AJZzBYkhbYqcrc0SJ247lRHAzNB0XPTYIK35KGV9AkAIL4VZl1DPDa2Zd7dLepVrgAyWDy8Wzsn0
NC7VHr8jFXFVlvYphaiIEKtNvKRDhBTbzE8G5xTo+lUxcGGjzqlVAvyN/e+dHYUpZda/XA4pVOUB
WjNAXPJigsWPlj11JmfCvF5LHMmOFGc+deMsHXub0pxVeZJX0Covy88Au281L+WVW6zzMH9abqh/
5NC3q708qyKZSDsfww5qjZo2lluWCh4VqEeGlHm1MUKcv/dJFkoCdF9BL+2D6O9PSGKVjsZgl43d
os8liOs+npjD+e0pFTAqYJNW/iYyOOW5jCQ6anlE0Kx/I+d/pFEwFI4ho6gRjDcQUTN3LsYesCy1
UjiLs/sLJ1P6iQtmWXnLCvNeYhJK6cqyXRP0CRjWQhSxvrX2QT14pnDIE9AqF6ba/j9b8Fd3YYD7
gbekdcQts7n8W1+7jN8ktwffRvUQRl8EnAB99oAl4alAbu6YHns+Lqh9o1C4ToM7K2dwUhEdUHk8
87tgObxlEbdwZn5qaUHE+B3yETZ40KmuO749yWk8cQOg+I8awugBSvuHsT8rvK5liOa/OQ/hqFUn
XLVFS4d9ATsqZqxYbR2XQ9UVkMAjKItBMAveI4xvI0BOoB1F26uU6bCQc28QU2pwgaQpO5VjKSC+
F16GhN5Chz+3sDUNqbQfWBHp580qCta0E2kYegfYjmyIhM+z2hLUH9BSi4rc6nqKGN3oOolk+JeP
rya+mzl69SgettBxzyeIkYWucViXRS3Djudg4MD6ni3r4JtYCqXPLW42l+GUbQr6h4+5WkDg/1M5
JynLhM6zb1mBjiDwRUcrHvygzbAmUz7IV/XLPm14I4RWwfM3A90Nejm6fWfmSnJwyWAiwSVHP/HH
G9dS0DmTeL/3Pd2GAi1OFK4bYlJSMVj4DThJSWwB13ZBeBGufFhEocBMensTzQsME0zTv3J9Iw75
TX3+kTjXhderbp3N4bEoaP6QFqsZWn/9VCxuqSdffWfLil86X9WMyh/HT+H/5LjVmCy4PBXKoLta
gW5lWGLCpS0FARcO0XbauGbYSjqNknCJK0pEVwhX4nXKonOCreXoayTe9vWKFJx1ALdKndJLgoOm
SwNauTw3sPwJf4ByVbGXdIHFveepfFfpWAZfXqwoE+hFydvdNWqpWYsRw5GYZD/VNqMC1AW0KGOy
k1x0TH0vq1goTXU95FP9+zXpiRAPGfLS+/bHx9JNP46mnctJ/bdSwPWapQs0+6LTvfJA31RvZFgn
aUo+N4ZPUoa8KFAe74xGdtRgq3hrs6TbGQEmg75Oolk+GKmy1WjHwjxZCBnS5trXI9PGA290PjD6
CQnJVuENOLeF6vSw6yqG/CP3SYIlaPjLA/Stp6Y2QYiOVmWhP42ceEmamfJRruhZUVN+RJND6tJc
rpEKIwlL6t6DnuMSzUUC+IYH+OtBEAW+DDMgUoabmz563SKVkkS+IN2Fx+m/ASLIBuilniGpD1WV
61BYDyWK50ooRp0or/1HC687MclRgnvu7wdSMTk8AQUcazPjQXG3vn9a6Wu+hQjEh1XW9+8CxhGB
y0HB6LkzmoiZz2lUbhlrzkL6Ts65PknS1rvWxbWWEgourewAs/mH3/WuIJ+QbUgTJlkV+TFV5tCl
hWwtHivfsruS5vRWF566YEx5k/t0bCzX+A9Z4J/LUreN7njF06eWMOC+e1G1PhTDd3fgonuj+hrL
VccXCsdo47HpRWZYDZ2LCWjbjayN3qeoScl/EqwzqGh/qdFZRyU1Q0J+SXlemOfg9LU0EaMg60iX
LX4owEclIl/yN8cKzGJnU66h2awLxZvMMPSOEj6izyscNr+vIiN1wEF+Ud5rS1rvLjZp8tyQ9wwq
dDmAFkEDUEU7ujSyC2aYWkVJs2oJ0LtCm3bdZuJLLxZoFbjwAvVyjF7H42NaxFhmSnYjyWbFAvpU
V5K9pQICbYnYC6uDx7JAmo88I86DPv9Dk1fjCm1DBDgPwTT6PP5/4daeNKvcRgzScbc55x5ON2Hu
pL9BJMPFIEw1eTUdrAPvwXX/8WuNUAJvEsxLkoeGmTBj33fmOyCUNUh887rIN/CvGqfaI/S1F3l+
dQGpZUELwBCs99dkjq44zY5gdP3VI33PkaXbxJJh77rma+k/JFZ+ORb+A0GaQvYALmnoVaJCpUR2
fMLanffN+nrAsEA/EYZnYKYMUjuFscIG6Wx9ccdIFSU9sMVNXbA/YAX6cQb3o2+5gqWJPyLk3eKv
pNFTPGEI7AK8wDXVi9kDw2MK/sqNJlL8lHXZjlVtty1vV5P44aLgJBpBRWdWGvI5rricCNpvnfWb
BkpSNEVEc/fK3pJUHReA6IFpRPPuYGo4A8a66tP91RKW7UqsjiY1cCFv3Kf46V47mEgLnioVBuzf
6N+HvHId+kME/lvZKHvvbcAuno8MJI1IaG5xNvXTdzApYZbvylD+GZOdigF88u08/toFHGTxSzSl
s82+RPbOUIxMNoxjDiwvv02UZxKlGzTUkZMg2jd+nw5t90g6aIdcu64XztlmcQQktTqfpXEkJQRu
WBFFc/2qgew7R1ttL8Rd0cM8e0JaRuzJDSvqkXiqN/5YLZ7nnhFilFBKtApZUXmIFU3LzuaZuybJ
+gEhM39F2yjVy9uSHgw5St5cn9CgU0ux+OZtMzzx6M4Q0G4nRvZvmMuJlK6133LM/dPqCXGBXhm4
fZvyshZZbHL7T6elHPk8rZXy8ttJTOcUjdbIP/DgdqZAIQkLgdenZzUYiiKPvuPUEUwecieHEN2s
N1Gw6trqMhntOF69zTCTNqQIixYtSXOHoCLVXUJor1RJp+F7t0G+K/YKwurrI8KWFuefstPUOwe0
zxISfbNTOV9OtHpuhVMghLyUgCrtD9bxQC4tMcGkM7IKjmJGcF+9s0/Iwi8bCxBO+jYWRSzoZteq
hdmq/r85bM7zCQrauJ/LqviK4ueHOVAy5DoFeKyE/gVE7hs8i3P/MlJA8G2VTVbmoFEe0vtP3m/P
ZiZ0oa9OCNQvrHfweeq2wOn1JLBnAEF87TOT2088ZMKoCf7btr+MiTC34YBLFG1/msKhnU9RKCIc
WrEi6vAXGozvOiWYpTWPI9OfkIYo4JcGONg/q+phN8wByh4306RGmbmcDyNIv8tKB0w/Dn/QDIKf
JQJVbJl5aitHPGuBZqbm20+ymTtgvZDlOH/HUuvy8KHrv9dnc8HNyUjGXkY3Sf0JtDC+7SeigStS
KfFmWxrJX23KgcBRlKewdGh2AzRfa5TFnO2sYPkX2NUPX5HRJ086S8BVtweFCjh3IzPZexkztFoG
59PfBu4lTAPe5O5jIUglTld0XotKSMtd63jAZ3ma7tRNWZlAm/Q/0/9xCAou7jmLkka7mMuXHwv/
JdWBMXzNNFPLwxHCQ4oLb7NFzcC54c17YZT75hOJEfozftLJ/P/8Mg4/jJIk7yKLp/9ebtxJaDY8
4YK4/jIMXFjhodp3p5Hx3cos9c6MZhDr8AhKuDzTjBeQzYx5e/u4wGGNL2AjSej810rtvBYy+7c1
9MVue7LmFVn0/qQxwkzL3nfcef6SuruZaMYBnlTykVJ3P5jbBJy1oMgYIYcEFthIQB3O2mAS13lF
GpyuWOV0P18Lvy28JfgQK9nE5FL3yyLzOlW9rbc1dEkl16K1+djWbTs2RIIWhmqITalDA131vSGY
pttRinDTxjeYEnPtZ/rC/6i/SU08pRefeXVzqaMAytx0sEuTWSPIlRK3rf0DkImfI13rtRFkB6l4
LKsYaKgJd0D8GpFKtN21nxCh7AUjptdQZpniAGp4HOYke3YLHMCeUn32fcUObDceOyhg5JwFlwSw
qVOJ+UxE7nS84s5Z2OwnPOiAHa1aSFOG9lucsMWJR8FN/CCyqJqMGYFx5j+ar5K+Ofc4mZzcvbVI
tNlD9zHAIY01j223tDs+afENpCjRxe62myJM6ykzt52xbcAh/5CtTxyQrFM4mZBIe4We2aHlPB7j
tIszBGYFLzZoOm/khSvwhoTUtAuBXX99z9WXO8dXo2fWee7XZCMvQpOLQhu4pnFZ3MjdBJzkSiUb
Ay5n/+KqCBlbdWOgLGbKSrodQ13rYcBQHzObwPCh5EDU9rQviaYFPDjd5fqceD8q7bLgqtqlyqbH
dATElnPsDHxnCXkB7A5groCs4e3CXZnsPfJsvigZQEaXaXllh1P3Vz6q/ug5JRnbUBzhkzYh7Wsb
YWxl4v9xdEzK1xMKOMbn1hrca1IHfU0JbxPjibqoLEmASZizfLE7fb5SiPF9WTdDNLQnJTLBUSak
8ien2TWbdbnAzRvU8JQR4J9Q6GvXPEYUvJxVUIWbVscTVhgTMXlc5vRepGlEenpFymEDiBZ+ylPh
hBvEfZTbqNjMukorCJMhUij4YY1emTVLpzpi+0ntCYJccgD99cUhIOeUjybGSJAyK1X2Nz6y450v
jSM69L9v97oOPOcgLzwgR4zMNmh4EUG/C+3Qifv5YNwhOEvLLWMEnsbwLLOT8xoT/rWgHA/RHys9
rcvqFoM8xXmFHV4dNATceMJg3KWyyrPifBaAHTGSnREwmwmHD/z4KgQLTVoHTCqG9JVTLUeAIKhi
D+xZpkNQ7Zovkw9bTl+2FI5rJa4C2Ec/AH/KrlSlxLi0OF0BIZYBI5qv2qbBBYL3F716xJEoB8Kf
48sDcldDIW7415BPOjQpyv3m8MK34qyQsYM2Am+DOU3Z/GGYTDeTc/+VF8hsM2CqQBBmFiaG8Sil
YD/tM5y3cdCfDbYvOodCrNmajawQPATjjmXIKz03kKo7AVMWq/LJs5WAfMB3jH8xvpYJQb+kLwKq
C+bA7yLZnPUj35AcX3CvBYCDOF8r4rDqPHoMtPGF1sPNVVcDlbBZK8IDy4SVcRL1cqilu2NRNaZi
ojzhv5N/sXSgnSZJ2P/eVU90IsBOOe51E0rEIP3eunB6k8wyiSToOeQynr9/WZu5R1lPQ6yEQFxp
MYls2tc0H2Jfcyc43E1s/fuXqM/2f7o1ZyMt1EzixwepRTMRbqiAeOeoO91PfkoSZ/bumkIOkD7w
pQU16jTSHQL//FMcye3aMwbZPvqFxMoaGPQvMBGMM9VbQo29hdASzTsaF/eto7TZ0GPwLwqP8acA
eMoQH7HRloz00Zmf8eNSDkBhSvWNG18oBT87zI1LPc2l+epRUSshMYZ4KvsjXw1BO7lt54uQBgCE
1O63jzKNbNPKWRD/dr8UQWBP780YpjBnnT3o8/3O28CNRBgwKPUo6lLVuhpQwEExekNKWbOaNd8J
zWnK6MmFT+VMubBtIJrYijsEE14SX9t/0PkvcsXsTsIX/kP7hkVPwREN5OiFTDtmnLwxvFRbfd8C
2AJRRoy5G2Pq9zn9Uvekf3iPakcC8YAJcqB1cVWuHjwhpA6Ynh4la5NeAefzIhngqUhDgnhSDPXl
1wvDJ4HBCe30u/4tT0x7ctOj00Y4XCxoSdTExmgOw/9HKYN6w2ZTk2vf07UP6uWZ3Jji8oh+CraY
AaZs7wTJkyWY4BD3NLkBEXbZlG6Kv65KjGbIvwsrBU4q2lNd5OuyQXc4wai/q7uRDui+blbDderJ
9cfN5LoL9cK1YRBhmx/vNTXoq11+/sUemjzqBZVYYXLbH7lLHGFax3gIBmi2Nqt8IyKLIBhqagsR
jX+E0MVHkC5IvYmaPOX7w7hnsgxJ2wD3bXdK3qqo2+jcidVdZ80GH7Nj4M5oKUiGhJkXcoeyNy13
o1rCJD7B5uNpP7X2SZJziNFVUitxrWgOAMIBaa7D6tfWOjdezgqgkCNXiZWuBKTBBSNoKunn0Dnu
StNONgDgJFYJTNH5XMF+4kiQjXTJSPlLlF8a0S6Az7Rkg7bLWQYPRc+I2eEJygc/TbQktLrr4vN5
oFBreQQrxJU4Y1/GpBdGU1kz3e8CoWWIR3vQlPQyx8jTAQl8ruMHOI9LvuC/M8ufHMDaXBZB8sMT
M9lMghw0BpUOZZmG4ZNP+50wo2TtH3UJuEcL7T/BcqSkTEmohwb9pSXPK1CTCW7nHEy/lKlDfAW3
6L5Y9+tzyzXfBm9p45gXoNgLqGaBTWE6Xcz2HMd+LKZwCISs4uHXgplSohV8fgTSUoGBGYSRGmhv
7W3ym2Zpsg73vNa1frTKvnig/PagX6FRWQvJrKqmImuYZnwfxtygpxiD8qEgHE6BCdxkNfFVX4+B
sFYZ9yHdGYlL3P+J+mXL4FWOmRY6U9YbNtMnP+JBUXICmPoh8aOswQXLiquGYpITCB0Ks+bAEvZi
32PcNafHCWhuOYNm75B3wQp5tuAiLXPljtxzj/z79eWJBkJy1euStFWP4HV6kyJevWXqmHRVGFf3
hCKcPx8Lc3IusmO3yIrxbFqwrHU8WQEwBuQNX9vry/LYtM7AZJpcmDz+sUQ451rz3NJOTD1/L6cM
eQM+7ZQWo+rCrxA+ShS5VuT1grqXYQvopTf0zswDFmEgedC2gcbkeNEGFVl9IDchjOsXdD6HDmFy
+CumsZf3H68ikAwjlFLp83jVVxeul2KnnYPe9aPzzhgWocULGSNbSklZo/+h8gs8l1JSkpNpM7vW
59uuJfz9hNt4bjkWFzI2MAtL6j9R1ufP56RdVC6qHP36f3ZuCH2k/Bf1c+P7nJUonIzqpM/Hb3HL
6nXcfOHhTkEs1uMPxR/5OVyoz2Y4vUJSO5AsX7SffbQ1MJA/NpBDdUOTCLYWDxGhrBz4VlOMEYil
Dt9R37GDZ2yzovXbAqEhpHS1TymWnKcIeld2L2kJuqdg3n4q4BR0HVN49og/c5zzSm42bJDp914d
2xYDExYSdgvV6nDc6QOzZO+G/XKA1ct9JZrfohs56FDPVhHDvr0YBBVqdnWtkNKr10vROP7PVNkP
FPahXWVVqC5o8ZnjtlJrQxO0oqjv4c699gYDPzaDlfXztgwiyveNnvIHR3sdHT8VmYjCrkTg/LVj
+HhvbghORfNCtiFQU+MyJLOvpfVO5up+EyQOCKSRZe5tXv4AzC7WMUpLIx7Mte9KokmhSw9KIDkD
yM4IWbqWO0hiPQjoOqjJgX/iQlM5WhqvpK5zdAoUXnxftsowB3PkOGbio5WHJA/2lPfDkZ3ItMFJ
RxMTN05ToOAYPpxisakca7qfCEX21rFgsei8mRfn/KQKucqhZmXCVSDpUder2Hkpl++4yd1pLFUB
ChB6oTlCn41NdK4sw++uHClQ9rgGfr+t33vkqs2ps6qTFXOR6k9qz7xiB4BVRcbGJGO8v91z3m6U
egRiEp7HZrWiT02kp/Fs5oO+nhlGA0lcMYxCdhJh/CuLopgD+jjcrK5NszXr93STI3oeLEFkx6nA
s7HeiDOP7J/43nzFg7QtQNjZORtZVekDx03aSxy5s3XSWYYeJd7ARwQvxK9WhYtZ8Y1MPj/ns2eF
hEo5kM7THNLtfBNqUk0cPBS7fFklmELeJployNOp2gHCGZhLnLea/wMaNgIphotkVzyvJVLElgDN
Pk+JO1Zhbd4Ym1Lgqj0AE3x4/4ovmwIZEGLPYekO3lzdMjiCXbDt3/tmVmXi7n5j6+SoXX2ILHGi
8ptZ7LEtE9lGRSfRdAcAqwUULe3+RWTZ9WsadvbQjWc9u6jrwtxWLNp9DW5p+LrU6Megar1g4oyX
mI/cd1gYYGn4R0QrFa56H4gguCe36KaQmQBSVeVz4vTsDJoC5tXUDPvvdJzJURAfmpAfTDyCFAGi
ULSsqh3hJkVDIiM6LU7N0x8Td0joWwAu4KSoYLwPW98upR2qlIDLUKyJRdNYpOxRtxFC0FhXz9qN
hI9FhidzwQwhLxv7UlRLY7YNGN6T2i/0oQ5JSdBwhA6pWY7u+uUsCd2Cu3rAB1XSs1o2WGDGMfxM
S9LEEEKUN0G9PMYAWADXL+vTI9L2dOkQ2oDbXvNOu8vxbmXeLPvhACczcpbePRXTmDXkon+drx1s
tobnRWHTKFglEl6q65qokiI5Tu8MC0zH0VchRpn9wCncOviO1afkPzKlg1U7086KY3E/9o6Iy3s6
ZAFdFCZptXhL1IES/L1UcgXFuyVtbKVi66ZOhMMiNlyzsYc2g13VULNhaNAepH+zSvhAhbyYKysO
n/3VUT38s0T4lb8V/myLRIjm/Cn9kBB4qkIBKbUyoVjAnaTgDKOPvY7bZ7n8OqAxb/6a69rvSrnO
ylzgLEBZmx20mfeu7D0wWlItD4qTIcQjDINBjzK4FNS4IiItXOFK5OczQYcLDo7s/+WzGmV1DZT+
nyNkCXZyMdPMcVbImY38dh+KhOT/pT4zLnOVKCz8NL+EpMJeUDHMmug8d/8XkLZCnn2LVaKv+JbJ
0hCAc7B15qe8rnYlFR3fSYz2DsS3Q/xtoyT3n9giz/NY7DZOwICwMBwTDH8pmzZH/CupCutUCJoE
V42e0hnnjT4AVIpUm59Bsg0po5xnU9/tnc8I4GbmyCatrkLZDv+TdVkuC0n4FKjw5gsmOv8SXe86
wv1fi/JXZfqPtUsZ2NYVK6Ny8GfVeRRCusezT/yqiFTWmpOLB5yLeCedCRlXbXMldyvR0JfoVbIE
LECqj3MFag0Fcl/wsgx9ah67t6/eX1Y/wntXnvKrev7mo2sEt3J/0pfQVb6FewdIkTnmYNt2BlG7
AqqYYvC5eiWj/D3c72NUHhmPRQlo6k97bPFOBcQzZv7qMFNlVbxBC0QIuW3JIipCXap3WqYe+8G0
gsAbEkXzGz5wszTHl8en/8UP8dEjImy442GCGy3N9RvE+ZusMTaVt1n2duFcyOyFq38z8e76rcMS
kdaUHWDlA8njvFXGbNgHgkgAPPHJya2I20T8o16FEca0yX5J6ggeG1amtoYr3eOAcT/r4jpiXp0n
m1ffOktSOurnvg51Se9ECQhEY/5UZWVjUAW4dNB+FC15btuy4bB4PnKSnGpb63jYLu+NGGgsQJ8m
Yig1o3H5F2mVlRFEZbi9FIXMHgGX7JfGQsVrGeJ7JAXXnhss5ogBPAKnVhizllfrMms0QVYU58xj
sbFosJSD677SdEyykg4WLG7YWZJ1OeoxVwipSwAwtio8YipO9au67R7L1xZ9ceYK7VQcivavMwx3
V4jRAbBP+H7vCnJgdj8wBhVT8x4bM0RZonY1vN0zxSqejFF+2T+UWli9ESB5UCYkopsDmGlMT28J
yQg/xNdJ/RncrMSLcziEQ6dCPRNi+iIT/HLgC/oMwOjpLaTHEsNwBLYwd2hZHyvDIbnKr7wbl5UA
arQUhAMrDMcxtOC8ai6p/wl+zRwfceW7LNvemB7u/nCKlTmDpJ+5cdXErwBcyaawNIT9QMHrIGbh
d/pd2unM2/wVSjp9neuruqJ4Q6cuIDyOaQ5gwvSF7ydOYOx+VokG0dxyWg+Wn16rujjr5bUDgeQs
h5s9I03+IBUVgegTUp0Ormzb6UlJ9P6LdLd7kJ14PUavUFkn5vcugTx7DkpTB6bxs6+CIZ66QYSd
6CMrckTlz7WxH7Dt/MoQG621pEOV2tnYSfHPvmMqAWQuJFx2DhLYuoShWOZLNX938VDkibTjpyCI
Ic9w3mHvtWYVAMtU8TN+WgDKLthLzgNwq7TXnYnoF6LTWxWwdXxlan6Bf03Gegg39kkbj1fS/JsE
iDbdmza0y6Jghr+drxM9X3zTpQMvSd8AkoB/QGac5GrVxkGHobY3sq+0MAniP/ole+ic8VgC6cxT
vd/6Nx9RQ3mDmYnKiDCiD1ws076Go6gGDF943FaT/rLsopX8IX6eH28sgasisAgu8YDBXCLMFgmE
Bb29YuCC3ENPnUIylKeoaehAEpKFJ5CXD50B5+ZnS7hvfOKIUSe0rK2NnvdBsOmzSnN8eTey5/3p
EI5klPENl4qUyjfGVVQ5pe4jrsEaQDjx6AW541OuMvUtvfmIh7y+ppzWEZVYE1q2W6QoRQ0tiA84
S7bXDf8M7N9+1C7U2EWbk68uS7rl/WmqERsJvuI5mda3yQiGluIsd6A+P5fTA9nq2C68wv2lZYuA
xqh4y6k/ghJmW8GYfrMBoA+2MLNqbCykukRuAZfJ6KP6chF83c69qNkj0thhz5V1NVV2MZi/vvt+
XqfLCssFQDgO3ik+uO/+0wf2hA1Z1zOLQKZEgzRSw7DLxeCvioXZSlatdJcekIXVjHswibdjQpIb
dZx154Y8VqlfCby1UDYAIl2ydLgmEZJfpE0TMj/Id5tfhSogYa7eI4ro5rSAiOAG2qyWKSdzBCL6
QwSjDRGCXTYXFf0QIjsMbapSINJsdPk/OdAjIlZxlznx+OANEDBUvSbwapGUergr4Dud60wtZa69
JkKHf4wAUL8Do90KoPNOhG1gjZqN3I+In2z+x2pVSHX62EJd5MpNrDY32Jq9F5VL/sOsXFIfaE8g
sjmKr8K8S6OMeBTYJnHwrIweLcLaOR/ziQxCd9auSBcyz6tbsfOuVM2YRogiSfEcjIhaHZcqQdHY
paAbTTF/HHLRYjpl5MSBVNutZCS5IlEL3YKWuyV94B+NGV7vVeQpjThInS+E6srERndNPdh6WhRn
6WgAq/yMtcR5gsfh5ZTmLThS9kIbvzXrHuUNGLyydkm8nCf9I4Wt/DLpwsiuh9PVKJQH8VJtkb4y
jUrZ8lYF63U9TCl1fuVvW0xImu4ckj63vbNbiI1hPK1Tfel/SqKzTpk/x5st+8f4t9tExPV8+Ayn
kSOKkan927RFGKZi+nvUr0upYDoWNyxPwzZ62cdmP3n3CwPbQ94DF8LhRzqUwQZthkdXft2LyJe7
9Bn0pBvbMJCWMQUKCCADlvp8WijEpOnXvegHQevuQWcuP36/G/PR018gRleGmTWgYI7NYUbcbE2D
MAMvl5Sw26pnB5hryYQNg12JVmkCSY2w1WhGOkP4CcKT7HZulZD6Jl3vA9tcFe8qWSjf04WBdvRA
0rYtzzaLDZR02os72b9Y/oCCWHtlIfsm+Zxif+m62qfa70kf377nfKj1h1xUNBUlMzY1cOYk0frE
ZGNocEVHk+sGQ0EkVYdMrsHxX8Rzh6HTrhymXJ9FGLTJgc93OAtnX3Ly7jrVqpqG8GUZCHk66yPk
N0JBkZv9UyRrw8jxInhZDv7G06sQYsPHXgDF9t1ZvN9boyQlxqT/jWSOdB/fwG2XB3xHm3JlElNm
NspiYYw/3QA+Akgsm5WNZZ73X+ozqGorkNpMAnRE5xzg8Dw5pDQ3Yli6TLBXlcNAVIxJUICTj2x9
6UeQJSGB1RI/HDV38dAt98wJZs/6w6ca0XOA6B/OKIokS+y2PL+dpRvdShQc6+fYrE2xxJkDhdkh
Y3km8UqawAAFjKNL4dlQ5ZoQzY3oQZGdU+4oiP7654qLueA5+pA/h5HOauR85dUFfzrQHtk8dKGf
4u2EORVqfdhH4YAD3X1UK2WTvgyuS0PQsyq/5scxRWNfmGUTH6EQljjWyyrMomwDltfeYOKM2SMn
eOGyqpSSNs5iCaAdb20RKh/9200djPxTQRVZgsATE5lPsUAJASeCvvU0U+KT71/mKkmHnUnZRIi4
1hrGeZQWuOeAdGKFLQPl/0Xa70cMDk1/nOXjLAlfqolaZgWmlHTbGrlAwsohkJszgg/MGAyTFoR5
CITLgFq/FW2NGVzGqDd0DfVcZMUcadd6SZOdnrtwjPNBY0K4NWezfxD454qEUl0q+VTOz3//WpqS
NWWTFeElaYnm2N0NcVHRF4TBKRJwQAwXs1ratig+k7xDUSKgaa15GuwDxL8TYZLrVNmKPCuF2102
jyCdjyQ9xPuKWkBuyKAKiER+JMCz0myQMgZ+7fE8Y192hDpzlA/rzUZQbx7FB4CaIzUk6rbNYEb6
aeESieJZbMuC7ncczJtMN8oeGlp+kANbmz1civfcd2rQ7P0DwVuiApngGU8mVzB8SEp2g+74dEO8
sqHffBux1aXwPI0t+2cuUlt3juaQyXuSTviXik8EEcAvBu3I0sL8R8WQpF6NvRxtC++yFZb50+zW
iNkbG7eCNO6Y4Paa+iONrRjDGTS6w+MtmwjuCXFY0JAOA8Jn3ZSGDC99BirR0ROER++0TiHH87xs
w5Y2ktyWoaB7/vbLr+OLefci22zeDgVN4MIFMbCvZhyrHtnX3C+RGQvGLWraxg21JJq45of06MrR
44p1/1uKKvsgN92ZJkCD90Uzov5EzLlKmo4zuWp7dzGML/1bN+EHDP45yXIdvO3rHjf8VsZZJlyM
O7Xj83aUHR+fSuyDjWvV91cvo0VJqSPYoNeRFethQcXN2OyVGIO2grHKn1lYJr4nA2/d8wf4C/vQ
4qSBRqeixcPOvFiW7mUcgq+ZXaxxG4iSjgwWyzsdnd94ixphtFWLw2amcx5Wb9D3qOizXQwM4SCh
+bn/ZMGkX+JDcUliQFzc7MId9Th+QIF4AKieENR9c1maVeLPwSL6AiPrdDQ22UXYwVkJOlLi688v
F9bnPb5IUITMoHsKv5zu94XkKVhi1rfkmyuhL6n4Eg5fDpgdeHQnkxjh+D2oDJFjKIUXMCamsNao
QIlNPvl6+0hMMjg5bDfwZa3UfgrtmUXAs23EFIvJq1xPW5MFHI1usltTLnxRz3gI5vE3EBFTrAju
ppXWl+SpVWV4MisxWK6KuNYRajiOmDUQOpQpURxrxxnzgn6q0CYzOH1h75rv+ihd1ampSL+M8YQ7
e11f4ZeVh6oFNJh60V4CDNKU89oP4n8qH3D0CLzN6+rDzP9jzrFAjrc7DjNq/fUW8WOEMFyGV+Ti
tdYwL9uAOyFrj1rxAbL0bF2BzQINqdi9wFhhopDFIHUa1df/L3Kj5cCm9s7eSGhKSQ4aD9Sr1B1z
Tt4lw+W3hle0/KNxtMORr+YDTkd+CtxTOyMGvPveGMikes3kmvITONLyrzhvT8xjOKjrk2uv3PBf
Mh5fxgmDuufBfpH+XfKBGPyTlN6iCTuuoG7eigm96ddBtY4lB2fwRSqX26ME3BtgeBj9nqv/9rmN
s98R0S9TtMwJHLWRwTaXkTRKV5xGaWjPpo0QrPGdVBCgFKrL0EZ91xeyVjLGVUBMUqmBAbhU9p1h
bYInteOHR9NCaEONk8zPYOxJhCdejLtHgXM5ymD5eHKSkl5t/HBx5ws0FFuZo171uz1Ey5hAgTme
stoyt5PJU6057VT0/V6iLQjqJgJ60YaGQ1QEnK3zr8iFH958w5tQ5rf7CMKuLJIgVH4RCPHpfTE0
5UTrxgNQMhuMZgbv55ROU6vRhzeARLK3Y5c1VgiFsDg7ITmdhD1XRFT2nYEoZlJLKAAO4ogwkeCa
8w1ORR5QA/alIT28oOhgumUj8P3vkNJVSYQnCTYCRG/ZvnP/Q8fZWsN2NevyUrCanpnMr93VkhwH
/c0WB0fgUxeDdkuwMRRqi8huZ8sUFY2AR53DHI9Iw1ifFNd1pctVaKwaX4ChwDEjBy6RdDczonIn
s/NvDgEXou5xLKspepy23zcjWl5telF3gMmGybhk6YbQefQe+5BNRxeff/Y7TbGEjjiZPG4/2GQH
3TEr/Glfd/t9y/C5yh8FYBzbEgw0PZyOKSK/Wygj/uD8teC5c0JgoDEX3YYsPYxNgQMVklDX1QQV
KckR5VEXmhJFd6bvb/L5sAZNONq+pnxf8pbg1g2/ir9c3vGOIYpFkY94cbkPWb489ZD2Cwq/ZllK
gK5hsA2RDBy7BJv62LQjYXNIEj/N6bhXh46DYkNk0PjnnbRmxtNapFAgEWoFMPAtB3IxCgMxOCMe
uuER+51YncgJYkE6hhwqM6i1H1fAFq9m/BBU8pUYIdQlchg0FjBKfn6W5VxqcyttiOLg2en6BMZ6
YlRykz9vKAb1uHb3+lvVIx3W3blSE8Liw1vAiaPThiA7QWOOHxARUyEjcGoGfHDX8Yc7Nv2EhMAl
/Vi6u8uBkpXtaiPlhiJzuXZPeJxXs+qIIwIlMWRSv+xBC0ZwYHTBTaF47LaVefywx36Yn8/07eAY
X+ZE4gAr9P2UcRim20iOazWaUGUh+dvw98mIrG3M6ygWjVv985pD4eNC0Smg4Er3XQUblJS1NmQP
okiuGaKPf6ltqez0i9BuVsMXs//9fbGvZvrRNCOqXYI1L+yv7G/Ke/KExBh0yd87eULZt4OmY+0n
CNW769JE6sLIcvBnrBKg64vRPAusMfCCMQWflK+vNPCGKK8ybi/rhQ607cfQuSMOo9bQ+leJbJ+h
JWD38EqTatY0N9BFkQ2PGi6t4W9qSyt+7TTzvg9ggDEUXoTKHJBC61OxTxq7Oq0GkCHSNjqY45a/
2daqv9P6oYCK6woNdZer2c93er8qdyVNQfC9JxEJ1/Y5+kPTePWoMnAJbqRi/TKERtOvx7W+vaIH
bq5PGzeSE1c+oug2iuXQHR+vcrqzKoFm9bw/NUOfDdeve5jx5C6cd0ooCVK8vBHImnP7bcLFLCEj
FmmouODPJo0hmbNERiCyI4rSticcjTzgd8TfxSlBq7S1jBLxjzO7xFSFdreN+C7YMcAUaTF8irC6
GYCRoJOsNCmqx4i9ACqo6AjKJQLtNevN9qjCYudMuE2mZfKwdb/0ZxqsBz6WJU90JRWqoGYEdXox
fTIZco0KVXGBX9QEfHRDDUKgC/wPBTNwj3BBQIi04BtR8qzMqMCXGZpCASArCMXjmP76G/8BxWYq
QTApNHSipUKWQv51j7rqgS9IyTNArPOEUVZy0MpGLRHAxvHj4Bk9CV4DCyI3FMT4tku6mCYXlMhV
H9dyXcRkVvksX/L11HPFxhALNciqHtZYBJuqLEf4Tehm2nwJwDAghBGSG+xsJ/r2GM/tsfJS/vwS
dT8tmWY+bDRJhjGQbtnaBWrvjm4/WOURsAVXSCJDgN3xgB7IKfyqhUjT0EBFKW38VAnPg7CTBFGI
c/SC2VCkaYZakSdKnNCuZXdqy5ZOQOJJ9yO2a461dnaAiXp3V3e4Vskzp3SA7tLs3ht/gq/nrgto
Szt8mVT2Fx0T1Szo4mrC9+w4XIC4dmDAc0Grcuy0Ad54YJulAXWUv2wYqoy2Me2cyHDpl4EAUUUI
Q43v+kkV21LvRtJoIHaiHEnfhZmmWo/tIMlchvnTrpfLt+1og1k61gMYxF4CprQ6VJu4ykl/MQUE
Yr8hv1pnUAykrB7Rmi6pKyX0lbNZKJX/giIIs8YXjflU33vR/8RGMLSK3cG1kmFFGHk2ySQ5ijS3
JTiw5HxYwcbhDTFIxuD4uyfwHnh29Up++iXPuFESwMo1/xV0bDl4UrU1qC9j0JVcaVYVyimK9pcu
F/xrpccWOhFlEKFFseYVS2u3rnK5VaYZWv35m+Lnj4xjkJy0DsMDN0fiRrN6aWxfRCESkgkX8oM9
1XqCqNGh8vGkO5KyCMQRF59Q+IQHo9wZAOqyKtdrsEv9wSwwQd2fJg+EZIr48JgLqKYcHt6FpN2/
AJtl5J0rUJMalZFqyyN5fljo11n6zLbZK+8o9zunZPmFRoPIgmnjkwQUhxXyAuYkgTKICuaRMbDh
ytp+Pzd+o4JIuCI9YQ7CLIW0O3YmYaplXJ6FuUX/iQEJEQohuPn+3SWb8DzCoS8OJ1eV1PJ4x53o
x4SesXpzQUlHnDdBow3Pjb2dTRS0/jWuNf2Hs+FU0dhVSIuBvwobN3kSwUpslp9jYequZRQVWnsi
vyFZcX8Gg1K7da7zm8cwecTwMONFYKwM2hHV9WtCvyxxE7g9Vx46154Gs6Mq/G0Q+ESIkgzppVEs
KXBxcRB2hBI4/1sGKrovo/UOcveI0Jb61T2A2lsYrGssLmHuzxcbTotVikr3IEh+WhYdTItkCgTt
rDbqvvSSfaW8nf2H2+7+rVHafHTCXqmBHaM/PTcOKTAtl7GjUE/+2ESRFz/DZcERnsI4yXcNLaOh
XbQ5izUjyT75H49cNIHbarxwA6NDZa43GnrO4aqUHUCp8H+rretwtDiJCFHI3hIoou2H0CYgd3Pl
YCFq0hmYA/QiRo8QwsbZLSU4S1ib+QiH1hYktG+3pgPQrgFFFcAtptNVNjZk+cQLo+L4tW0NklH6
fagpX5vecis4hetCC4yOkXGBzjdSEFQl1m9PFRjHqfSQBAN+tSlFLC5Jg5crwwzEkpMVLiN2LVjF
X7vBUXivaHhgWG8WKHReOfhhA/LI8cdca/R91EnQoWU9U53FJrwnFVJx7iDkSjgtUtM/dN1Tr/X4
WujgOXOQNN+tWGcgSfFDeikdG2cmDo2T1xaitpbNN7EkYcVUkVkgLKHdd7fwArdhgmtrTvL4J/Hl
V9yyWUDYnXq+KG9dnucK2Y2z2PfOU75a+/mll8fqm34aJSbcFdPx0mywVpZOJv94d9FCMbCIWEcd
J77n3HiZOTp+lydqhJ2VMe2ROtA8hqjvIIca/pSlu9+AUcPj/49ZqzYHaCfL6lNz05zUKWtPCk41
Ye6vDp9QUDv+bG/K05Enp/lsj7TkeoSwJ0o85B/8p6vWPGl4WCGnJOWJW+pvkwv4NWg0uDYx4Q19
NiFdp94lQbH3G9fEQkvMqKH2RFYi1vvqoVOXeFkcwkqUTwlVGD7RKR2akPKHOKPXBBlJMoakMSmZ
5iXUM8dWwIDtsaaW/LbPLvKlROtqNf4vpo/RP9axMI3DkKAkdAiqRvwDqQGZShZWTkqsZpvcgefn
PUhHfjQ+RcekAFBOhswWyds0OFvuqym/9VfVmNN6fKX3ykcTPYl0MpWIV6TtQrHm+qNlFCfpRv2l
kKNdjFq0znM2hcgnnI9f02P/ZC9QJV75KvMobTchGOkCteBMjCTnyK6OaTtIzrKpnWcVhdgeE+T/
W9rvg0Bmaj5KmLzdU1Lx4uLcmg2sHPkd9H8AyJBN12OeMrDnaaJt3S9GCmBmn3CORx6UDjQGBLwU
GQJXwWQ9a4uox1Qzd1zzuCVnZvUHoj9vM6b69xj/pu4QZpM5/mFFSIIHl8W1i0U3FYR3Z8hrWOCa
2upweNr2f6xYXfGCkiRU7DjZHQchzAWuvpN2vdmWDw/UylqVnZsE8fGooz6t8EHC45lY9sBlul0N
bqoakiWwZWeKsuyZZGjaH6ELzwGeYZgTFYy79T+6DQ/w0Unl+4ov7CS56PNcV5LhBYxHuSbd4PkU
cKS2DQD44A+crdegU/rTrTS4zgW+9X9R49EX4yPnhjVKwCP75ob4O70mg8fw2rKOv0p+wDGmYJ7q
qqOhm58+lhHBsuVzbfeh/kYuHQc7LAzimJNBBXUin2NLG3ETfZAENPElyj+IFPGmL0Us7+8RPX1K
oClhbnPlFYcxDDzoIy5xTDco2tgot6JlpJTzJTKs3DwNznjaVmWZQUiqIehphacMDCEWO2ij/FrF
nOj/jjLwaNjJlW+RSETuGmlmZVKb3SdNhHF5hTFJ8TNBNT9A1P2LbzHhiNns7t9aqCJ9+MsfXUZj
ZgSvM1Nkp8QilsIJ0j7UtQnIZn5RmKTc0OUb5lkvRkBXOHXy2JcVqTU488AaohIQRLY1/xxkgjkk
0YSFs/iZ3oJZgPewdJgzCMi53yHpR6975FlFq4dkNdHayyBSXGvedgqDF2zCcBxFOFj8/AkjXjEu
4/twLjG3sVEtUoaPqy+hmAPFi4g1XfV4jOivytAW+am7JPBL7lL3rd6giVJ5katmwq78e+nZA7HO
mtk+HKKybVOu7KLaHeixtFyxWUe1JExljjY4gKEk+xVbSVAp/ua4lN8+YH2h/PXKyrt70IbzATyh
nNZbaaH7SxLsLSkYYP3pnrBYmx+ORSu4svtwxqnr/wOYSqtxmSO2f67+L1xKXoHmol3H/jJesNw0
f3QCEN5RhaUt3jHF6FpcAj5KkXeEAunM86V7UUfW4zpE0rK6XKEQNBcmWpRV9PYUN1fLUqFzeYN0
mupg1F50newS8KlWAh8y9lCC+neOleBPgWU8g5eTF06zqWjmRCnvz1HM4cQYsk5gRit2S+iLtDif
gJI0om60kRf/Ruln1d8vIDjAQN5eY0jd/dT9HyRTkbSGbha45plkRVEFHUH3RTMjMK4SGc226oZc
hWWGPp+jCQ0om9rJwCmg6mF++NH6zYWqT/BLaPclRdzQNYESWvV0nkDDh5iYw75I3PjlmoTImIJ2
03U0S1nOjAn/jYJGxRibWz8D0yuvz1x0MArVsdJ+qR8SLzvTsbxKo9wDJuaa48g37KaQ+XfaEtRD
sxWG1K9rK0rPZyYwUOloZ3h+5YY63EoRUJC/P/x5EoY0ydl4njGmNL8yTfCJWBvMdp0ycf6kfFg4
YJQhNLQ7GNpujes6hZbdU4eOzH54rXd4TVoB+dEnxXlOpKZDRawqRNM4Vvg0s1DJLzmxwFtLYEKI
T6WD/A7Zq8UO5HlLRKMWbbpa/6DCT5dISmC9x7LoAhqZ/8zr04W62y/AetkjtNvoaRlTGhu9FFnk
wIs5phbcMxu0YwTE4HIpCiSjYjRFP5icDVL4VVAqG1jOxgEFQEgzKsj3qjJsnBk1WqVCxEAt/x1a
n2ze0oHxIHscEfmfSqi/cYD6CFPQhtW4mxISLD7nIcuBsuJd+CmGFUdySvK9MaDaGH55VRLPA4cZ
b969tTqFjnbkCKAkfM+SzE74KJyW5ifwJfAUzDb89oIWq7fOxPQcpEs3xy07IIjFdyNLidJZS58G
tb9UshuxPL2dAbtLzAgQsCkyHkf0Xc/d1bptE5LBoOdrrGX2XX+2XJ0Ws0XUFg48yDhF23MKncui
eaDGqzWp7hJvaXphUiB0apf+DRUtaw/aMcXBB/kFT7l5djfm0eU4aRsP5cV9PaJwHXpsvWR0SzB7
FGXfYiIDqVAcfmnTIdKbwotjnyZ68EKNh7QpnM/VTfhrhNHr5oTCRoiMDbQXtuzi/Ojr4nzzdCdf
dNKRMphPsq6Zdlgvj4Y3RW0ctApQ6EIDZPLDisPIuXxurcWMAHpTaU7kmnF3swzP7N4GUe9CiBph
Ofk6zXyOfMsutDErjEJGibZRQ/oCn0u+VNcgq1VTSJSp1Xqc22Ng1z9RP3+W4gvBteA9CLyfNdQ5
pBRB3z09OENT56/8S/RTlJpl2o0xQ8YMR+Yx8OAX58h+39h+wkzgci5Raxw4j5oMPNkOqGahDJ1O
cXxclRNFrot5jL93MTQvhhB7/aLqhfnKxqz4hUrsxoJ0hDr+LtTxHU8mjDz+wLhpPaBzc/0wkb9y
Vy+otMO/eiNSAQ1NdFBSweSjYUQ1/XbEgEtRQoy7LPzV6VdgI9JH/8T03B9EpNcQwq2bUEQNy3sf
dlaIhx2Xzeg7JrCoUTt4FSJJga7tFuD3uTMrzMaPxONS1MkjBonuUFBarM7wQjd1EE8sgm1rgYM5
NBa+Y0dNUaUVGjwv1WebjXw1LdioRabxju1wbJsYVgxhOMQUa4EGp1qaGMqPnsSSE0UUFbAWMCeb
nc53lxgfSR/nODudGQMbXcL/iBNxEYMcCKnQfNPhi6myRAJLP2d4k3IUZ6Dnpyr0zBTVCT5tLEd1
03kIWnzdxIp/BR/5sia3lF3tKKzOX4l+IpOBEV2mI2VHmoKvs6ROvdHHLfHe95nndMQxtCBUtbPQ
IlH+jHjUSr/cxnCtDuze/sopkYZ5veqV3sO/i/Pgx8Cl/2cKJC4o1kDMRQcY6TWzoa+tdJwMHunb
jmejT+wfRUhCv1o/ZvJu84xzSi+fnQ7pZ5icDXbXtyEImtVyb7TVX9sqs/vOFcXk3nt7DmuqxS8w
n7snajbG9rlC2nTXVzCawnFnHEIjBZSiug+4Yq15VOzzfdrnh877OYaqfw4K9TtFSdQAV+5gB0eh
g65kYC6uzYr1a67HQEirDIkNELYm1CQw8FgzSne49T+LX0ph+Xxbc/dHLx6bYR+yMg3B4kZ79R0U
a7c633sCdgEb8fUeaCsY5CgnZ1+bqSwZgBxyXIlgi5GnfcZLj2qro69t/15SokTNy+svyTP14hYa
ehsfTc16AYIVjpdT3Rgu08DBetNl0ZhWFtGklrmghJprROPQHAUpd2tLvyL+2ZDKZ2nyOe8ZLn6O
40jcv3qwgdQAbSXiWqEY8nY2gS7HnBcHm85dh0Jl+cOM3/YjD3+AzTZiHLZPvxve08CB4cQ8gc3l
QJBr7AtSmhemMKf6suiq/XJ7wV3pnGZhs1INZViHvs2/3O9QjuRVRM5UfHWU7OmH0UoIDu1Qt5D/
vdeXlccNc/Pcuxjgr4Xp+PGMdDPelEV6m+SXnFyPet9sC1nbmKafTLZ1otj4XBpB6IVzreHqT99/
qXzBTDJqU6YAhr/cgW0/ox9EbEie/RdZ3vY/qYBmPfHGANcDiM44jiL/4iEios9N5VWbaHR5ZDym
B2/WdZkOCEz7Ex66RtRlM9FnwaESc6DAnkkDYFR4/EH8Nx01eEVmvSiS1UdVgUtdQapDMQyA5PnY
OoyFEThjA9pLqDEzT/uO/bEFA6GRkZ/bKPaFotJy2WHJtFcanZihs2gUd6GRCipBM/2RtX1X27eS
OowUVWyFknqdtVCMwvK7GorTY2i0doLEZl2R0LfA2IMA4Fa8yjT0WmU+7m3x0t/P/MAYLHiN26Uu
mcTeS4UGtIKiW/gJMtPDsgG2n9OajSxxOl6F1DeJyPZKdAvYcgLnsGiVp1hHS5NAIjeExSTElJag
PP7ge4SV2+kMEDGPguNuK3/Qg0gqdNtP4fwv+19JiseSDSiFMcrMjp4SpzmAH3wMKycxljft+MTL
b707/pNvI/6HL9n77NtVKI7FOUuMwdvaWZQYegAM62Lh9ubnyLKFvrpOs0eYiCDzzrRPIN/1cdLa
KYAGfb91E1t0w2JbSRY/lCmTk58/XDCI5mjt22fiqkw2exaAlZEk6nBnMLHWXlkHm0wMcbwr36vY
X52jQ+HLkWmr6qhPKH6tVtxTBZIHXjY8mzwJJtYK0WOtHKGk5QDjZbpf2Pa4E6RJZh/XSxotF5Zh
GyjefE5u80aRupSsyWOyvBHRi484b7pRKtN/GH34bBQLqGBBcqOCAz0O0yii2HrOJ9opYmV5wl5f
T0q5XO1ceiDNbZkUz27amXzEhCiEjvsB2Dpz0SQEHom+Lz3dHQuf7e80TnsdCXi0aZ0b08cbU/f6
nPX1mP3d48y71pnpohA1YfOWpXygcYu6SPawMKElr+uHYhfiddteRoL+kNUp8mPAMWJGo9JpkEc3
5E72jfESlPvRcUt0Tk1xMop8PFubMcNXKzItBXavLfwmevVN+VcROsC+q27w1NxH72J429jI14O8
3j44z4jaF4Wacfnl1mBdT6hf0hH1Nd+zXpysrkLEi3Kd6WutXOGSe7U6WZ7XZis5nTD+4tv+u9tN
eMah8sXi305Gqu/JXEwO3+gwqTySB2OKI+hZcI7ki+Yx0dPHXnjv0Wdd8tomSnplwe1cApbW+OTp
yN7gvamM9F1Jf0y6mSmZ39B0Va+07gEdXrVDqkzfN2vhBv5EamRYqmc/5dxYKLV2nj0bmkkwuMZA
wvpBE7WNBUCDYC/AbrQWBo/eq9LsrhT+aoY2bVdu97dOTo8AbARqhALeiOLQEkHanv5/HENg02R4
6zKg03nOqK7uXIX9dVW2yHme13DNAVEJHof9+TbaVrd7xPTwbSpqcy5Clvqkn1Q9mb4u+iLU/Uiw
7tQyoo7xvQ3a57/uT/W528oYkIRlTVRdHJ4dPTnHg4h8ZKANiwPLyr8MHXP4oKSRz3WrZYI4Jbyw
WR9Y+7JfLXnApYM4UY7J6PmPclhLxDI/ZUI7J0J0hQtwcsO9zWiGzHIsuxk6yGeDP3bKVwhvrO7a
pvkg66JJom3rtQsoSPVxdyPwETlkZ2P7+kv1y4+p3iyOlquR679dGwcc5nNB4Uq8qMBGeDkGGsKJ
aO3H0gAlZSao2jLHVZnGnw5QmWi9d3/jKgzrtL0a8smyv215Ay+Kyrm5aruCZWk1R69hwizY85EI
Coid9HEMqqRnTZ7ibEhHZXiEQtyfmJWPZsLnr7twEuGYW0yPzFUyK2RhboG0IBEhwCyeJtBmlGNN
Rwm80Zr2wj8LEmsCSmPlkmOKdOi1JZVxwGT10RuJwfbF4ovoFhLQYbK3y/iKiLb7nyQGCsWZ4Nz+
HRZ2OHkmKvsZ211eRZFrHtv8ejnIR1W7UxzPdqRxD7CMrbdwdLacR5u6f7qOr5WWOXnHLvn/sxx6
+edDFxdYf75DJO76E8g9D0OAFJa+lqYoor4itmKgrKflKQ7pHZ4e3MhNnvrucg7mad33TCYqqcMH
6H728E7sjH7KAfArH8r06X6ZCbTQ9vG32bfF+RmlJ2gVU5dkC6SAiirRZyL4JkP0S/0MTrvEZHi1
Qq8qoC++C7HB84QVbqiNpsFTMs393vjwFEC1mBiYoDVaxdLtMLlS8DxfcMV2027Df6J1mf1zkNsI
2qKcXqV++7CTnuazUbI1efET5jtAkmnky5p1/49R7lautZQalbRQ8/0jzD2aVIjlUPb3zUZqt8JR
RpVJ7NX3DIU9Gc2CIJ1UGVLS2RccFBsvcKhFZw04ILLyoyqcvkDLKklVN5n+86Gru0pbYmK4oOrD
6uV7QMWat3EX50aZuwkE4NxoO7y+nFkEnnWva2u2cpgpdMCFtVaku4tRHadVMfgbGPrPW2e/oLyD
77Lo0wlROJvg3FQHndThFjzIIaRvyui9ujv3DNTIQzgPjp5qtrnWYx0USXRDwwvetMH5kxEHvhc6
dRB7kO3GWrCsj/NKQk+64laKdZwX2jsDCT2EP8AuHGK50LOEMCzSJdblM0FKh7vMyZwLIJfZE+2k
Ty5iaRBaKg5UOOQs55FnINJoGNlJY7SEIq98SVVPtJ+RKOa1B4p/VKpgBxUIfxxiZWz9lRWvRru2
tN2+YXT1erRT/VmOtCoAb4xo+fWOA17tXhQoSfF6/80Ez8WIellHgJWgReI7jBn37gV38sY6mSln
tS+eI4i5ML7zjRrJqto4IK7nfPYELbnZyPKj4+9wKBrlPo90GiaKbrSoyYo63WeHqyNgfp0y1b9p
k1OlHY1gU1bWqxW11upr4Cr7I4oXsNeXYWq7ynY13LrM9rAQ9FVvnaI9+SGcXPkfCPOtYcBvOUjz
JMIxOnhykMkcrJ8eSpnyonwu7WaXpmfCTMQP4urCxtH0mSRkRGHI08P0qUu8PYjIhiWUsuxOSJCe
XumFvZmZDVaKaZ2/qDcNGJKIHZIADeuTxO/UOzevgQIiI9kKjYAi6/6zMBL49OloU/nLhbEzzEQu
FLOlx0poAyP7NsOElJpo+OYkWVEIW7j37IcLG2ZMNywRinq4I8LQ8/4NHA/9S84zrOQdyWA/mQpT
jiIdh65OSi6PepZzgacBMT6nnNcdeCVz4NxrdH2xRm+rm7X+bMTizZMatDoy4mDlcQaHeGjpI2iB
wyWMScEZ6W4Rel3+EBrtvfOvnI3YHd6qfZ7KvrXeQwEU+ciitdV571Rx2GjcSTNw8hHyoN7Rd3A9
/dH2XkY5DGO4xJ3B4TLUeDvKClzBuXtSbfRucthQNB9EKEoXOb7xCUBDjMy5EXXSSU4fOYEA9upQ
GNMb38HWbi1W/jckGwAzTNT31pVHL64FwsNcvYTKwB0LSMVP27/kT5P5L0Y8d/vNtVURJ4gtjJwt
OpCPdBcsEbUxd0/62RAPL9RZGrVHhUoveE8KOM9O+H4N6t+j69VMHmvtxe0Dd2AWXo+q/wPMe3ZD
oN8baiSwxVgX4IJ2ZQ91xxBzyy5C8h2alwgw2pnMWy4XuOaAZ1Ds4F3kYZW8oQqo5Ybt5jC0pTLc
t6SF4ybQ2eAVMwYbrl3bC1hrAgElaszwkD9gWb7ShttnrBMJbo7GM+/Eri+kOuA/qgAl0oJMDIOg
r8zsAhu1Z4yN1t2V/2b4eAaRh99xpGg2cUctUIoVQNgR9RcH036JqAXGVppx3CYAjwcYGvVVLTMA
YQMVNRBt9ujH171SjRqdrXXebQ84S889ii+wqgzbNjHzSRxFyPeplBZgaBusReOn+WCH3Yhdanfh
VTdricKVyOgmrxIPGuBiE026b9D5U+8HsANaUZ5WmOYVlvca6XDetJnIXQnq6quO2/cTKd/hnoIZ
eoyQ/E3VndpuWrEfwxXJs8uPf1AFw+cnhZ9KdwtEVlENMMIs4oGYDsvzwEFOD6bDL8xWGtlO90lB
XAMRipHHFpkUWADG2J56/arBe55LiXPInqzuiVjsiXSQIdHNskwSVF8j8zloLGtxYjNOpnWDmyrR
cixt4B3ahla5b6iz/GaSsZO0cOvpVwvxl2SbBx8qGudduxMXPnyb9Nx4LBSHWb+5eS7speaE2bIX
57iGXwND09SAKKNuoKgk4fnQvJnk6CMtgjpMoQcKuAaq2N/UvNHOgLxiMZfD+iOhGJj656xe+cQx
Ug2RWa4/8vKwRihIbddsxFg5Js3gRFJy+vuJ4e4T/vi4Y+bVaqnUTc9+Yv3FbKNtxrWl9QLj+wBU
FKaSvzVuNasRRnnTHdgXAgrF5s2Nb4Gf4JBt0z3LyQH0+IpfSiN9d2x5RVJkqJ698Xs46ScyIDKQ
pTv7gAeHj7tIK3SGXZkvw9Enc/Ngb06r1J4rZ98Wmm0idU+TwykIreLjLbrjxfyuKpeDS7pkxEhy
hbJNa+G8nL77LAiHRcn6/J8211Qaegp4sxvWjJzM3xzPT+roNTL3sF/DI2l4I8Q1FnWWMPO3nkjy
uhKaZ24l+jphTzOMQefEA5YI81/ZfMy9aoVpMq47yg5HO62K+WyNXKzmoXUTx/j3yLsILMi98Qks
uOdXbIIrIKu+X4Xt9IWECaICujL03+Af2AISNc/JtXEBRKBt/FEpXnFon/XCg33qNSL7ux5k+y7x
FoVUv7p9j8JlvFQRwIsIAkOHqBjM/+4RsBauoIxc+EZjipENI/h2YLEpKX3isTHAzlF4woK93tCg
bw8IosM7khyWo7jxugvoKRx1L8futywKGgV7LJCFiqOhtiD9HMmE6cgi6TnE/szSLsqtVCxsnp6z
IzotEVDJJtIg5tpcR5+iJrXhJ9q9PyJE4b9wIPpWUQ/Gu0u6bR+j9fnv04muHuWC8YwiD7Jrddr2
LImuKs0Dz9sIe9wLDoa4L0gSrgcUT2BlGVGVkyieSg7g4Mc+T+A4c4Qa85Ua/bCSTeYjQG/Fczua
9PhoiveZFP6L6o06T43KiRAZbFcwnlr7ictg4Ne+d/aC2w+XcUfduq9Lh53amkC0eHIXHwj6Dy7F
gt8JQ0q52zzy8VvMvbNzXK+o1OCbVkC7w1zpI7sTf9dmujBxXXmSKaWawcjfUig9YKswGlOvt1uA
a1JAUcS1tAB+dW/CJBWNIXwkC+zckAYB6/FMmKLqoqo5zcEKL3r6jP5DS/kiqhMjBcIRbsFi3Kf9
SfYZu/SuxC+7RHnmM5ujqKwXNvINL5t91aVoErRDQIehrIt+zMRtExzik6KEY/11spXtn9znmH1h
2EElJyg4ZQjTTtTL/dCEH63WCH6ydMES2xC1xnEPSHwksfJ8Fg7DGOadhCMbndj+mbkil7FM+TKN
SgkE7D5tAA7esAjVjHVsPr/EzEIvnfRYsgKG0kpRLukZikCUBeCmGxk5NyBrIiO/fpdVjDmeaJ/9
wDUwCKLRWR52ZYsUGBzWvTv7A+XvNdHWCUFvHlZswcWYozbgF8wY+LiszXwRrx4LV8gmNuqeuYgF
Y9vcd9UImrPvejkmpkIUKumr3cMOlkU5nzcvaet9nLa8mrdKdZtEYwMazxRMdBMaMAYM6ZKvEcqe
S21hXZJslzKyg8re/HMSE02qgWAYLKHAjAgz4rSRSjI3QhQqEozfzwESwidYZyIbggxrcijxtfWu
+QJdfUjVFVN2MjYnW7RVoJn0xLKzt0rRbYY5s09bgINHQABzcQRjX2OIR6iLPEvkS1Fkddea9dn9
p3Zj9J/edvbQa4z4wIB+yd/f38oIdLZ2Rnmsa9ImnyXxV4bdPP9xQWDU3fBxr9VUwtBol9KoJ1zl
T5Rws98SbsnTvHVe9PQZQbrHusvIzvUqeol4eLMps4mgvgrTUSC8+BQKObatcFXZNlMmNediK7uL
+Ro6BgcDciapAmFxCQ5wxJalOVyIh2jsyzs6jEFJeNbj/AZwmSNsp7bt9UKl9Y/DvjHSbyR/vQW9
TpnvGF67x6MBb5W6W7oREEfPVLnOSX7zDRolfcwT7PhJaU24Z2vK50oQun6/9IeZGE7RYIpMv0rS
OdU2sKKnEm1Z+/JpSoyXXQDvCyzubeoU38MaDkMFDgzJNeBkW5ZfXP4I84skLkooad4aRK7UWNVQ
cKNR47iVJSaczAjhmb+LFN4k3yp3nTC44/XopBiH2lo/mziryJUi80tRnEUCr/4/y8AbqketlaHA
sThamyK/m2GJneyAGENCpOiNFP2o5TfKQf5ilM+rramkDWAhjKEZTv2JzhRYjxJKwJsSLe4Z7EX4
GywLGZGewtrD3Lev2Gr0u98HI5Y1zkKA9N2yPY7U69+D5jiJw+64ZeJr2iTXdjQCJjSOcd254Txa
sIiEyqKW76pwGgLk9zBnechV3UNtGKw1fhnGhmX9X+p7dDiI55GQI1z8OOiW1JZbNmz8IRx47ECA
mzzUZraPbhCxQWvB7HsNoG0/ByQ9YjyQdZs9/gp32pHbVK1n1ydqUr9JyauvQKmyPns39xBrhgBX
VNSYXAlX2DEhcBX9tTXmMFmirbxAB3g7VXGO049Uu5uSLfOmqloiWMAX3xseqG7roHAJGDxxRzBE
5CODlUM9rC5VBjV0UHTSR05BQMSD/Tq7nLioWWthrwxL3LRU0tLaADEwEblmQ0ISzNmxRgj6p07L
fdL6k1/OFcxFdNtei83YX1rXwiKCLSx0IjCpqNnZR++FGDf4LAy3EBLbaRMSjTBVdDf8424MIP0t
cbWKqjcrzAALYUqozwLcexSzz4kbO5eM563YqaUUJ6qjjp2SF7AUwZB9BmxiOZuxZsp1hZu10/aq
eMdgIucdsag/sas6jPkMovozc0aA3Hyhu2PqLQTR5XIvL3kNCoZN7m5GdqFVI3cl9V/1zy+kpJ2f
YaMuvmerB3Ha9Tb8opGp8KTzmp2vMIdVQh00p4/0IxGUfKfNP8VLNkxY5kXvMm8+75/c0kcU8Qb7
509CaDb0yuFo/cg94syUwbQf7N+dUdn4qerktD1jsZTAjpvQhD/kF3ZFBZzFsFtIQOba1I6dKNlb
ZyENKyL5l5rE8hXaEkZKcy7QD4m3ETLnE3aUxgoHhBfswRz/17mJCuz6rY5jASP1w5SQM1wbHlCC
NI8P5te+vZpt5x5jickqXX+dJr0pXVqm1gOqHs0H5b7bZNbCPIuWfdjE1sI13O8bXH+2Ns0fFGf2
4j8/6wsOAlTH8PK/PiTBhS+zjX1qN9kRAmDV1IP98E4URpgbKLg9YkDqPxDpG4S9WKnc4RtVGweu
x+kMyOQWF9N/7hu/CEWUahlnAHg1kIwmGMmSTI8ZpkqsLzem4eP8cF+oGfxjAQ+5DEwEdsVrvfXr
iDYfTgjvH5jhzQkhKuHa5es5ExxtKxXSqbVaPdvvPfj18gmv++hX99UABTX0zOUo2sVv7m05m+c+
jQqKHT2QXv6lUc47jvNx+jWblyOOEpn+8zBQ5hAlciwUAxeRJ1OEVwckCthL61zd7oWyU9Ak8NLp
CjVdwVNdVenY+ORUZ+ye3Za2AWPZs624s0oQvzrQ/pFAOETqIlI0dsgO6FaW0fbI68EikxYu0nkp
3YErwG2PvYREKj18SuKVNVJUgtHu1HO+7KSr31DdiPTfFyCMjWDr7Hal8K2/FgYLhR/xKUKnzDKh
VdNRX5z/SQuMiDqPsp0tyuHfEs06nIorYROPJ2KEx2ZPj1PZe9k6u/QGXedgdqflNg9uaOl2apHx
WNstczqhXLLNMTJY25/eJ4CnwxVv6MbjSyGkY6IT0t/MDX4BnVByXoki65VHl4wOWsRnRvpMXObk
EBaeLHYtkBrZrtIOk5N9oKzwJZSscTXvTgKyYs/9i+6ZLA0qP0Kv4QoxyZyzoxv+QHXQi4t23Q9t
AUmh0XDwVDIeWy+6GuNktarKIUAmFsONfs6HrpmP3v4f7HYCdSTYWJOW0nG7viUqHBRi2Nk0UffJ
81vzY+ZVJDxLfWVVoWjKCkz3KHzRCGoyU/UYvpFBL17SRKw1qOBELsVUEJJhsxj7r/WHs5i/k9KU
TyrM+yiv9jaIMt3Gcs+Fydp6DJalkN8q4bBsxS+NR6BlMNRSbHC+ai8EQSidGudHR3HRkbsC9YGL
gZVP1se92o8S/EzBq86dvsgnT9lHLOuP2vaxVEtJq/ptBGJ1gP9X0IBcKhqQW85AshXAu0Pwesrf
7H3GLRg+eXgLtnXv+0Yh7FItppvHcOkHLUkDJJuKe+Ex+8N6NMUJVvY2nI7Y9ZpMOYW/akimJRHk
v/JGHZ7G0FmNYWXefTWFO6H0EG2bPabylwpZlEFV2grZUOgtSe16nySHVJNNc8eqGfLnhh40X2H8
if54zp94Zz+WpPlqJMFtM9GmkyHZEvjVkaxe7xWQqiKbFlhdYJ23fxaCOA/KbO2/hjqhlGOSN0Lo
bAtYy+JklT5a19Eg/umhvcYTjicOfUSBGddWNPlL7iDneZGxfgX5DDYLBC6f0/fjuuPUkn0z6Ywm
Am77yRIaZRYxwXnflj8M4LMqrM5GwZKurz3QXTWYPX16CPuzMLGyBqgtqiEGKmZXCglpWb1XzGQH
9zK8EshSHf9s+OqXRA4VD3zs9qLR6vBujdjKglPeY1c4CEYlzw8f0ewuvRheRwT5RX4G9ncTALwi
uLw3auJ18BvOEbVe5G14t5zOQl53mWiXha+M+gMS1OjvYLLq1NfiQpif2q87lFA8zMNbGErPvuF2
3tbSCyLv8N1Flf0Z5UqVjtGgTfuSICOvJDbvoWOzKrbGfruOUk0YPoJTpEP7e3/RAL0I3KGLUA3s
y6j9JcneyrAsuac2AgicGxRaHus4W8QespNUx0iTPFx7hX41+dZYIJu6QYsuagmECgndEz63Zhtg
MxVRr6i5hyq59ihHEcKGJmMu44iue2g0iicDn458WRIdkP16NiOh46IaodJP/YWrgQbMVCZo6KyM
ZsJ9MW2H8lAlYp+suuQJuuA6FjcUwz4tYxsODyBbJSv27xE3ZtyZDZFH+7XmzM2ORTLFFq4Yt36n
s9k/dzUja50QVXR68PeAKwTsFxy4pyfJaTxmBwc41gWTUd0KamfmAdSrvNUx1P1xB2mWmB+0/JuA
+6bm4igvyuxguamGCifjYi0p14T3ZVSEbVx28sVJQON/NLXufsUYspC+pbXHzhVaUEaZDH2d2bND
n0dxWXB7JIo4/IRCVTmLr7rUD0zJIOwc7J09T+FoMwuqVhRgxwWIZSsqyXt3mRSzjecfTPN2yVYB
+AwQ4Itvnej/N/XkcR7L3S8PvQ9377xkNGXdvhhLPwd6zO3jhOYNYDb9eVaYI1hitpVocXLVXgGu
r7Icz5Awb342jxmzy3A3DDyV3zswJsCdykeFF5xbYfZJZAB3zN0jKX4er9E2m6jD5xaXMkLF74Pn
FoH3lO5TqrHl26+Y6sJXS5SzwffjbRMOQY1V6iAKat0GVEdmn59SRssS2ENWMvfpGsilxbveUXIV
bFFYLSkT8ZczOcTRH0utNzj65ORvVtGDzvyAE0XSCRlRn9yOT7n/h4QRdisofVYBBG8JdHQ709vR
2NaNqruhi/mDCH1k5beBtsxHQCAGQitZBWTjKigQEq51ttVaMLAzBBHpypnZNCbztOCg6tu36sPb
FCgSGKMXy1m0LvZWRlqyleELhSPN/wmXc2PjN5rNPy1Pe4Wen0MdbmucXmKuZ62EAEZJEzEnISLn
rT5bTdn152kPoHteOyeWZIfdCyrZZI/fnxC2O5h3zZyMYueF8Fq/I+XEC1gj6ayNv+Ysq+VKgYsI
I9V0loiY5U/jJQfRfbBDxPQXj5zW+HCfsWVRlzDhFd1x5cvfzR10NbmMIDGZ5D6xBz8sRals/1Ut
LBY4VpT4HV10+0TfgXb8fNkfGUG8HseF9sdkwjSUdT3t2OGnyrwJzB9f4HmjAm1gdpn5h6V/PB+F
s+IhDs8CyowB/myVFECMcWbYKo9Avo93Z2C8WdVwwanZTVB11ptVrwrhxNfcpYvj3UHYCxle2A88
QItYwsjiipURX+EPDYANvWckzNLQ/eLdB4tO57i2wVaNMwfiEgxv0QFY28tdc9uy4DF5tyIqoDr/
jdTkJrvj/fgZf7CY1yC/8OpxZaiZIFVFRr6b51pI+oA6dbqFPCYuFfOpnXpunel0XA0jNG4SLOvw
qDd1tWJa/Bw90ejZaqGIW2TLJGG5MG7/du9MM17OgDvhf0n2st8WObd2XVvO6wOBHm/grMnl/XAj
+QXDRuurT8J75H8k8XImP1DhsX+xi70Pp/TL0lJwEeRG4qDgaTxofL9hxxPTp9nh4jWuGXDLLGV+
/05Vmn6Axx0q4USuWb+HuQzcpa1LjKl7d9caKafh+kzKXee0weZYsmc9X111HpJNZ64R30cluNld
DRU32Owz15MOkZkqqrm45wVoJe7hJi85mNMO7IPSjGYQN2licAoGDW/IcydLUukqz0SHtqcMOBQo
71lEzTsbjzPnxY2+JBRuJ012WTtgEYssyq5xdHd6AGuicjosxwA+USQ1lQvRvbWywSeUHdGFSALs
EULClJXIIN+OR36BVjzTkin5DekESVP07Aue6HxT62eAlKsxaJA7458csMxdyyTfGo8zIPax2J3M
65rcjHyvuf4pQO/p29DXo5jqDUjPjcbcWV24ZehTUZWgFtAGRwDh69fEUccpkxby9wD0J0sGoqIV
p6lC3Cbpb/Wbrhp+l76rVA1sw+3oDHmj5K6SIHw+BbSr3+RYj77QTXwFzgKOdzaXinB27QnPbn24
NVlxzYo3lrHwOWOinazHCCKpzJ31PTviKrwqvonPeiMqBd22Rfw9mRNAgTtKVNmf5xAKqIpOWAUw
b4ot+pz13lRXj9E07kVPYP8TpzACYeLufWTQ+steCSh6rJR3FH6ywJRThwVj8RD258B5pcoPcaRP
Mf9q8RqgoJr7pht523PqR8tmIsBAWGmZaXZi+PJrF80Oa9E04zoEg81K8Tw+0p/9yeXh8JDvTxpg
Cyfoe5ZhJeKUW2UtxsKFwew7epkdFMzxJWlIkMCSyi/afCN/uPqmjtceYnKbU2Slw+Z2u4vybwQh
78N7A7HG9TU8eN78EB51Dm/bQjqTlqT2fBdrMgVgT+6KHOfepdL2pywmJDSLJOWjAPhzWpCrl7Jc
RYlOMKRe3wHbhANqKZxmv92jLZgTlEyvCfF/yDqGM4CXihKGO7PeJm9VKkeXQWwVQrKYTqborRsZ
ykdx8CQKJnIXRRqtFvtsGk6pptfpvjbinSsm7+aWWP4tbBULrO6GFzuwLlYsYte506tMpIbBZdIN
sDgIVkiYkMsO+24JSNK7ljGZYnrBj5oeI0JAlAw2mR0hxJKWNrqr/pry3/wN62x+33UhFZrddCXr
kBOAvWOTYNEmD1zjHTOxE5Roa0USrfi+sRUrzFLj9HX65wpjkC9cTdO3dqoL639ii39ehquraTAs
V011oZBOI8FKEh/jG7XDpQGMaAyQ4kAj3gD+0JjT1anV5apTN8C2p4yNdT8oa/DESPxpz9VR//lu
kB8ed1d6smx7W09ozZXLol3kZoYUxgpyy2+NTC0CfSdRfNxVc5wdzqUPcBi6IDi0JhNwqqhidGOo
9QYO7RpL3upsolCLCXxVKYQ33objv3VgiJrJxdVlstAU5tbYC8V/FBS/79DxMlVfZZEMVrAy+DBV
zbq/Tl6bHGs17Tmk4/AkuG41iDfiyxWPXwmlZXoD2dHuYYrPA2GrNfeIJ1eQYTie0b028j95nbi7
Vj6iWjq0j3uGB8miJxHC9pqMojGGcdd7ys9Beb36Pg2QfDd3lsuwmJFMdWAXIRTLCoPcmgcs3eSd
w62bQhSSYpsqzoFPFpn4RfAyVURQ6mG+8O11xuLP0391XrQ96yr7u0ZcKHUYuwKSzu7kF0glEbXY
SMapwJ4839iPOw4bUnLmFGye3DkurNc0Nc3OklXqmn3HeSe+yXISiyF3LnjIvzL4Gv6f4WcS4orL
2B47sFMWtQPOjTDUEJFTcce3YQsVLwdBF2cc/fHdFpP4yzpfvr2XlkeYlAgR/wPZ48rHxeoUQMWj
zonQlqngDZiEmhT1gOoIXT5Xn1gcq6CC1Si458i4bTRXifX4t1BfHQbjJax1snwHUogfPcBC2Nkd
Y+OOJA+xFP6iNDJhX4l8uT/GBIhmxleC/D0l8n7l/VxhlLxRV7Bk8gflIPUbbts6AXNpjwMTu8Op
7jFfnysj4AuNAXC4YwMNDeXYzI89sMTuqND6PPO1m1Tp5rzY9ZA4ACZP88P7H5M07iHo9DZ7KN7i
Hc0Cbv8kRxIg0+2oIyeymWM68gzdWIRIBEgNO/BWCedLmvk3YnOf5xwH5vjmQhlBDJKoiZBA56WG
Z0GT7ZsnZvfN/Y/l7B/UO0QC7Y0zcU5wcohBkDi4RuGzxdv6wJjpDxSqxh1gI2doyx3GJFStX91W
h72TWGWgrS0QBlHYp/IA/6+ICnxqVba6urBbrbdUG8wWcYkh7GNZG55wsCpze9NiovxymWN3t0aZ
4IuLCJCfnoapQWxbthIlq2E5tzD3Vdf37vX1qMxuhFXrP5tSkPV8M+3ANx/SNTloXS3y+VzzqXXm
k/oVQcoFoNj4+Y2WhAp5sgQiX9ajMCzB0FAvigkLCFJYqni+zgL4QmPIaH0Pc0rgICaiEVxA7d8p
bK+yWYRPesvDAljvYETPexoEu00llqaiEhM3baXyBzetHtgoIEEbkqrPy+CD09cEzizhByhDLLXY
z4cxhaOsIdfpCFeBqudtty6vEHyLuxZtjNShGPvjo301mx94T49Q6N5N5TIvobgzUK/3GltMPgwG
lTTKkxtFpCvW7d685frHK/v+539kXb6PW+pCNDA5JDaRH+rHlwWzD/kb+yWRLgVC1Zw12NoysLDy
rV6L4f4DDM/Jcyva+ir23zF+yTX3iyCUJ+wGwEg70seZkcEfxDJAp/y2D8LqS50bapAw5+x0TgL8
OUTdOnzXmipa8az6iIEPxno1gzwu7B9sfzYU3A9yitrSWLp/1RUTfzTyV0PTWcy9LqwWhNJQTpXJ
Yy4g/CCwO3n9vnIXqFZj/hNubz3TYaqk3BX3qHK4+ogQars5MofJZnW9hZUvl7o1DJyLv2pQpZ3G
fx3A5lWOUFpDEfJmseT5Feczr9jMaSsMu3Ng8hFExppojU7bAEuOP4tAMwtRD2vCI6G2dkX4A7vh
Ow54FXJBiscwLESrioA77JR6ux4Yt8V1E6apkjAbEdiF+itJ0qKk0e6OZuhoqLkXZcS3T4T8uT4n
/RozXxx8FqvfXSUMP/Kufq5PPyZI0sxhXDq3z/i+2BstpJlrh99PTTICjCQiGLMqrgZkkUU+ESLv
I3DiUzlD6c+ibSlyKxU7gS5rq0vjoOYHoZ7z8bQdpI8UeouLNurYlXDaI9rFZy7jQDX+LKegbLiT
hzxjFX+/X3Sv0ZI8RNP3Kkq13ajenSgBxVnJA7c/F3tiR8Oyp7KzqQg+wta7uovDVs7U0FYFnau3
jnVqf3ztq26gGboh+mcrP5hAp8SCTGOVZ6NTKnBb4ALZ5E40508oGPU/40tRJS+aAZSuV3skAaH5
UR9CXjL+iUBhXTSjMQKJeISFk4MtPDyon4qFjOeN+jV6o7IvWYL5LdO9t6WSxAXjoqEHeGHh0Ggh
RueoIRlfxLWMG8EizBAEHdStCaNOR5SVy2qSp0O1I6E9oMdeYniIyn0IB8TdstVsm89EpRAcm4Xw
bEdc6ynxjNYdVgWVEifMaG/HwrIe0UwHS29kgCSadES7ywrNQ8S2YA5KusQpol1gMAeBhpOk7EDx
ThJqEopuY0snFG6qtUd1aZxiSFIXQ/i7Bje+TuzQfj2V/9to6FHFSsJON2SAaxYH/ungYDA8RqoQ
Q/VDcjlZma1JtUvnpsg5cZ6JfEGxxnuIr83I2eV++I+sCjx9YQbUwjgrYMR5x+m3m4f+vJ7PwTLD
blVEQZB2k7+zhBobpc49ucEN9FL8OTyLTLPVPgd75KyOP+Pztg1ZKudGvQmJhbvgnGNVIBbEsQ2U
oZfLxMZPbQS9zKY9hY11UHlTIaq3Ws7yim41WsLRmReEkkRXGwjyRJYrmqrR7fNaWu4AM2s2y8S1
UDT2JGrKKczuraA1Sx7qVi+35or+qiu7Wdvn/o1vGwaep2BKWnSTYpTOWQ4uZXKops22248rmTus
rqGqn6aKoo5rqq79OcnkRqNDH4ULDF1Xr34UrbGnsmOQroQmfuIr7d7tCWXg21Eq9x2YKtAul6cZ
2K+W9MQsfE19Q8IABLSGt+W8GWKp5oOUKQuekaWLOtiFdP3ClLgXzqlRshkOwAfSge7gJ5hP5ccV
rIQMUxz5iiZvmB0N+DynhnkLvscmFEWac+ztef6ZYiHKl3IyZqnztEThPmhtLIQEp4SCpdhDzuwY
IjRTwZHrquJi2zIaWVpihCk+q8BI9NzGtaejSSn9UrB0SOkbJje5CJYljDpGQkk62r/LTlP2StvZ
26uEFVC+F7JIiR0/lKZ/MlQYPNcLkWhDEHAyhXmQMGwRiQcbRKz3YC91eCVq3nPqEufIhse0inNA
AOUcnomeuiJCO4ib2P8bMXT+Q+W2JmC1OjTH9ezSn9VwDq5bDnra/8SxSeWSIJyiZtWgHD/nHthO
XSpLJCM0hoJCaFOLXaB0MDzotkst0D3YRRx0Lo3xNZD2Vdn3pS8KuEknZg9pyvQrdvbky9hBaeXL
3bE2Hea7CCP89jhj47slfrGb79fM/5oZ4NUklcE20OXO0Ui/Lv6Glr5SuyF2c2HZs/p6GB6/LNER
zRKfSUG2uRsBPqxZF/SAT2/BBG7f88tnvd/3Arxslq8YmtWNJWx7lqMrufY3TRxQbyqcyCNTld1D
ED/3h5Xjt+Kvf7jGcwOnaFaIiUmtctLgOyS5l6NVod4WhHqRfE5nLYuhcDkSvP7v/KmrEohmk7Q3
uHy9rfa4llZFGmGjbM3dTxvxpanQsFOmYftALShYvQXBbHMVUUhAEOi2wLkJAE1y88fchVcC2JE7
h9OxliDsjsZ1TeiENJJ4Tj1bFzyPiiuG+P0Q9H7DIVkpsHzf7NZrkp9IJkelyT8nobcM37lmBnaS
hCrIfVLzYGVfXzQNVLwhUGz7D6Hoj0+AqjjBo0ZBsqLe0njM8EU47okNpI5HNeN8zado+YbkH6uP
0zmi75eeHg1mtEaOEDx7qEd1udSVoSyJqX1skz/oinHifMYKoRyavv0C6yDvIet2Rilft9zk8h3f
DxyqhE78cqao4hfBjvng8URj1ESRNY+9sEjvqyOagde8WCGUgUFJjKq4m/2kZ1aoTbsNWrF7kH+t
WsZhTv73JmximoWzDTCKMwoppId3eHvwTchz/IGybJlgvwpDhchDd/GS43F0/3ydfHckRhdiYSYC
sh/ud5BCgBnGBfJI/6xwt0HF02ravwHsAyLdK+PDlmcmJoT2m0jR6XqQ0NRB/3NNDdaRbyuky12B
FrAZv8TYEHjqrpXgkzdDMeAJbbfIanZuQodpQxShMMlwNU9FCn6kcBg+73OtJiCcA4fOz1/x33Jw
h7k9YbiI2rV3abR5hKRrR/LF2em6EVOrgv7PLxM1tuwUKNFpTggpFIY+MyWejuN2BwHHdszWwkcC
VCky9MhhJH/ntHJWElpFXEQ2qVfhThNZI3PJZ/1FrCZePtJD/8l8x2dp1t0g5aAP4WHZj+XI3ek9
ykVqnxzf+5IPqZPEdPu2M2btvGidpPuyGBb2v6Alq4BbGXqUCVkHAeZwmeVHVdXOKps/I6Cukzlr
FKCQt8e6ALpgz0Bn10YOalPCNxp5X3ahFEH1EPHwfk3Nvzboi0D3vU3Knl5BZAB/Zk6fQ2zrHLHX
5VTwkW/PHlAEzX/iB7XkEwOdvKkW0aqv9bPqa/9+IXhBt4ZDSX3N+z2Eb8rL0ZSOFO1hKDzqVc/I
17SZFnfirpsgHvk9pKxC2nb7/tPm0EHSfRH30gC067t2nVIyhNVHOYj0ZZkkgIqlP+ubYbDzn8pt
7JC7eS8Je6ZnP8fSytrViXHTLCQydXwX6M3gx3r0ITUdXjfJyIN+rEJNTmWNSWaZzchgzdrHdidk
XLF26J+ei5+QVyS/7pdpvS5a8B5nOgRainOUcpWAElYF3i/Y6D0WAztCX9SP6j3xXnvWIUDfXeur
+RiQJAPqheMQFJhsiwsZJz7iaPznUgWYE1Rxtl31+ZU8+smdmhf2FHSpwaQDgs2pK7lpnJeC2WC5
ysk3T85vnWQhAZrrOPC6pc1ao3XeQhpj7eR+7zG4cmHrmEnogDp0N1+Jk5FXiX1v+2RMZcW/bIw7
kHfiP+5Y5tUPfLeJo8X4AJ3LUODtJ9PR6tWkgj0BjCwUmXg2HyeBJ5XymO6SXjTdZ7TPhR6PB3cf
7m3uHj/a/vMKGVd8A0zy3B3FsDWIFoPVpWBfh8aVeJSkBT1ny+bbzYtDFnZVvCURAcX+Rlht1Trb
SxCmM7a8ra9+xhjN5i0sHcRSH2xSlipi6yHd5oMaXguBn8W6oKSREwSMcfiFgB00aILU513xnCLh
k+l3ahDySMdDux8Ie07hKPiftxanU95/jweVKfPbCEZS1epzF7MMUHG6FSKx9FZGtCeHnLKYFcsW
HV/BCsszN8gS82JfZP7DI1r+GVvvfroBxTAl1gCIdRzSPKrB/RdRI6VRBp1ELO48g0zC6+WWYBku
m0uPmSJUWSWo9DPQmMLdOwvZVV3QamckRHbp458YxaumAIEG3FfiUWvYaxqpSxsfVRPB7kmxB/m5
XUhOwHFlh7n7dJvrmaYyAKt39h6NK+8XbjDOItUCClH/Tg1nHiNvTz8VsxltKql51V1ZqiFIY2EV
GaehzzLYQwFCxZVeEEH9lFzUZU6vU7CIlL5hNiviCg44ZDyq4CGx+sH1ObEmPkefOyV1lcyrIik/
UsvSmohWBek51ixm6mpBEvhgjOcrVsTi8aV9+YAOZe9HvpObGk8DuOjgGm2VHDN+S0iKQI5OTJ40
CP7zXaFX/LhhH1B9FsVpBifyo6Kb+kaIxtSWUEymHmu0m2zQO+VZ/VA1tWPeetfG+s+MgpLeU3YK
NoeNr3y9jn2vPoSGaphmcsSnL2D3aAkehNS6e0ERkbxAwye0OyCAAKEUnThuMM5TxUck8Q7MECFh
BSP+rc8xUjBCDrLP6QD/rkdIOaUkubrV+tkrM8Lh/2fGyoz4blyVRK5cq9FUtD33Fx/4jZvk6nVo
fJFVmWv+a7+eglqt/E4IFErMsytxXOQ+3eGepdzgJIFxTGUWLKeYGVQ+k8N8aO1IXnfHBf4enVar
Nnq6ldv+sIYfc/sf6qyuEXD3SJnDU5NMSLxH0T7UaAWY/WU14ZhfHNXyguQL14M6aBJMu7LzF7Y6
lVkZTwfqxCTkfrcEoUdh0ER5FkRlBN7JXdFogRLPCXfWbPuhX/tNYhQJ0GloGmOCryL3ami3zGAB
ILaz2fKl1mHoYA2l3TqAF3EmFiwDHEjAgcCq+PsuHMmZfl/WmpcnIzMN8Ppgak1UKwwib3RHUy59
is8hqkfXx93PC9Fk+GaisvLQ7MNNveipdURbP1kVSE8WZRkzsEDfk7OcKBLagYTMaFGSQ1tqI9ku
7Mlg2elgL82yD+PIMJWJHehmEs+q3VIMf0Tgs3OcgnAhEJfI8zSoXilcj/DREnZ/D6rVz4Kr2BY9
UeYn3+XU0w5N9HebwBuflEQ3jFcBuMDcosiAgxiwqM8VQWDQ8WV4geD+aYhZwiHkkCaPXn3pYXBx
2lOfDH5JVn5UknGOFf0k+9EyfOnfugVbsa4Hkg8tQfO73M098XZqIvmdOfrdEbSoWhF7zbo13nJK
2qQxrjenohpepl13S1ah+c4yltb+pipgzVRP35etz8UFWdODnyJFC/AsNhKDH1rjsMMobCjFoPCW
9BP90/HucGoNTMKV0bRF7oNP9q0y8CaYWFZWW2McnoymmizTSljjx8uso2ZvVzKAZaS8f9VPK1g+
GLbdoyJcgM3ialZ5l0vt9ywUrUbqD/HDURjjSw67rURLGxMrVE9jfQr/kf1d2o4AULMc6WMZFXbd
YznsOer/p7EIIEayo0Tn+79q7tL0TEhwvDmjAp5xuXqvDnJEzAK0VXmgtbxc/XPZXexhNErnItTI
bysORHMMdp5FuJRWRYZLpkVnOUFhtvIRa0dRxi8eJ8XTwDc5xhEfBRQvtZjWWQpW+dgAPxwVF913
GK4V/1HO25ede+61ZP6PHOVEkrMmCojSjBrEiE7pWpwxr4xs82e50ilpc2w2BYvHbFT7O0O4iTvq
NEFdg/Wlvp5Fx8fe1e7r6VOeDt32EqZsp1eWyYtvWgUghVoYSZicinOGtAqzGuMdjY30yrgot0Ro
FI8ilzdtwWs3FVn9JCecz9B1Aiisqjk0OVujiBEnvmXiM+yR7rpW1irx32tM6G6QiXItb8l6if95
iUX3ChzqAwjDwPEC26yqyO6q+Bwf71AhB8VZuDLnUQvlGpQjC73dpeac4ndEcdyRln4WzecjGq0Y
j8wqBz+gDjvgReCSCy0M+7sYfarTzRapgkdaNRwaDDCnJ8nOH5N2I6x1AmLHC5Hk91ZYtvO8yX8N
E3mLxRmoaVRXSR+moMhe84rH2gF+OZ+2VWGiXeQ0muMF72gHOEX3fjCIo/zGqPJBmMyWJQsQu8pz
P+ZyusXwTgIVUjyYtgvye6sdgfAdYG9IgF6aVIkwEtm2GjZglwdNlRARBYXSVB3seAI9nZgMACuA
JsMk5nd9+GzniMf/GkABRCeSi1aA7yVQ4waMlst5geVcuOqQP2wtbuks3prll0DlHJhBbeZ27ZtV
bCFtZUjc5KH2RL7HUKidBYzBG0g+BokP4+uwGLm2Kny5sLhp7zYGkvDcjdDn9KV3Hk/lyEQ55JNg
iSOl7sTuymBr/GfCnUCzcHcVbQ8x2r6lkzTaUMHu4v+27QdzscF5uoQ1ruxxgUOr16bD++8mO3Ao
qk335m9rh90JChWQ7scwfssI2mtYtrr4F5dcwJILlyCDCcSqkxB9Yyi053yt+Upjk9tbilCO71D1
ilSa7ko0jv0UzWood71dICi8Ka1V5IMfB3fZyfnwyM1JnvhXshN1WtOkZQqTUpjorYKrWCK2hajt
h0AM1jJTxLYqoI3MMDWxQm0Nh3zSU+xvuvM8f4c0m79ij10huqNZ3xkoa4okQqwlGi0Yo/Ba3QPK
2/ANc5PuHeA7nlCuBJIQwuEcxNuWhOhBXU5EMKN4uX8sYcI0bN/8nr8Rf6n9vSic0nBTJOEX69oS
bprxciKoNtGE9IaTdJ0q1SKl81WB1Sawim/gfL+WKD2m+XIWm0YocoUGZ7DnHGT3m4GI6dpyq/bZ
w2rlRNnX4+lrtvAkfGirriEqU/8cH7x+WHqVP1RmIb04O/q7zEkVAjPhCeeba4oK0MMs1HKU5nFu
OSFVwJuOpfN1xrbQDCKenptKFbg72cVZxe/lq1SWJJ4VG5sQ0hoF7SK7ZBaxs5HroBqmzkuIYO9w
kd9xq8/PgHp44B/PL0PP7l6tadgDpJQCu6DhIx9IxP9c1SruX53n9zXDF4JteErkIJwOjNu/ifJn
X3vWBEtVVY+WzlwJx0h9yehQhZg5eGr2iTi5nErn+hkf2TA8zE8QoGcL5gQRkOgC/OYLS/XT00O8
vV5pPgTr1DHNQsmBARbCvkzv6qT2op2agvubRmILXrwjvdDU58dPM0WtnvRX5ZihfPyKReA5EO8Z
dZXP7Xs4ktY+rL8OcMaolj4BOupNlMZV/8yGVXaov8pjRuvYJKzIDjIwA7raAw4LZw5r2aIye7TB
Nv+Moa0OwKLAOmuO1Q1EBg7EmwMzw43CRcBExxNRLjtQH0U4nRycyc0SjTMormdoXcMwfC6AQnPe
aTyEp86+GPjXl3bWqO/kHsRIf3bD2hB53kIh32lzXuWEqciPXbigwRqhE3cGCVncWJJOKkaEjrB+
wIxZwDVVSAPwlOLwRSNv2ALumgRvyGys2RR+AW/Z6hXe7Sre2dRdsO+E/SDhwjl7knDtzcDmgszE
Ub9WEy7Jh5ODIOTVIQWSBFLGj/jK4UgTwIfYSdX4uMfxQB/YKjLXrdRKHrUWxh2ZpPOKOUKtD6K1
ewh/Dpndiv+BRyrUeQKGtwl/6bvddGSTqbsm9s5emp3nRggMRwFrzonUarNKKyskYsyAM5nQkWQz
vS5niqPEr7POnuYJDnxQyfKPwY+2Bm61ksF6GJU9A4UOyno5O75cwyvCU95RuyI+NtOvLzGSuKXm
4T5eDAOPdr9PhTR2s2bOHdCu1oOo/DMCbfxuGaXmI4kxY5YyVxiulHG+LMFBuhz8yJBGZRx7top9
6xByIpZKCpKc0SGV1QlGrhU4BrFJF9kfDhCUIOt2zFCrgYahPX+aTfF1qJv9vkn+R2rFB9lVqQO7
oCB8/j2f8f0Yr0m01W2y87TP7UFv9OuNvhONDGIFUCjnY6KhPqRAiS6h6JUPGUos9DgYnQnpKdiZ
B+NsEQ8FKX+in/RzBfnnE0nr95u6v8OthRBCy7MdUdH5rBuV9K+SgBDywCVRmIy/aAYxm4ORXech
cLour5vW/4iRRMQS2D+IuB0sx9DCZpEvgGU/m4cSR/5Od4JuTPDnbGW3bbHDLHJnlu+dh0dbUOXm
7qEKWXF12viKBATMZyEf4/K5piyJ2/HL9JOcwIvVuqSmRGBXti+/weYSu5wBIW8dP+HBjFE9UMKL
nYiYYID7hj3c5HX4RZOvUhBS8xhsAqdPFGGnRfIpuBZQqk+6UuK9LASikn8Zj63dPzOdoAbbY+ZM
G1smkA3maKUG9eP46mRZv4j/gQ3bgLqiK1lGhQRphWrIN5JYzCb0A2ckeZMgVcZlWacAVIP8DOin
enb1oWs/+zH2KdEVkr5zYItT2vJhiXqei0d3Jvg1Bp5tBQgHAef4GkSANjSEmmjB7T+227po4jmK
3yra9wcZxRtGqUUAEBWqA4x0+ZJ2BTZQRCvfvFunzM+XDhDGZi+sbrLndTPT70nn6lA6CptdJ/je
oB2OE0NgkgnFADw+UGVwm6NVcMpXUl0xaoancMljVwlnrFov9NzqK9Tx/b0or4hkHrP9WiNtg2Pk
Xee3PLzOEP8gj/xxT9hgWbqaEKUHPT+kWP35W5ZrbLWJUZk8Opr/k3//wWCs7XmVfbLh6kn1g7RN
wAvB2A/E90AC+4d1f/ytasBUNb9vcxD95ZA2B1tz0F9xbYC5X67Bf7/ZafSC/kv6JzQehdlgBScm
CwDTCWVFdiQC/I2adSdKfy4ugPnnIQfVDHBTBDtV6KaAFl0YIAtDqqqkfwGonR9RPTGCMawA4gwL
wLXsHrQIhvQmFP4tfLSkwuekiYHu8o1pwgACcyLHr2yFgIMbKlTJRmvTfimxO95XnxzfdngESt4D
Ue/kEoW6uNwmmznsuEki0/lvRO6bKtwTfv4r+uTEaGKDhbwdUww7pQplNvdLOg95w3TdyvhqNbCs
C2sXBR7f2nZq4uPK0DLxwZPbQGRoyTZrXb7U0qmE6MnGv/hOC5uqx3qd2NKHQZGGhsW12efGV8J1
FUYyxiw9EvfeqWScrjEwOXLIUPVF1xUeJF0jVsWkY/9Z0RfLZJtPEI6WYnCW19+bZ+YlOS+JJw6T
x7eOEKoCAGUdAH4vk6DiOC7FCssuFqbL8AXjkfiRhnPDvArDfTcnF9bQp7e8oWTZjI1zQl9YJ8kN
pomhS0avjBvpMRjwEMJ/Qb6FSBlYRDVRlZxj9wMRCgKQ1gepIKgDCRlY7c8LPlTz2qGSm5gNaBMh
FtzLs+sqFeGV+dUCKXmweTv5f119aKErJpVFo4b3KpNRR/W/CkaGMgnC7mZU2m17oSuPid5LU/iN
KlGxnTaNZE8GQSh2+ucmLZVkl6rcr+Lz+fsfQZtXn1Npcy8JNX7sxU7LjmGHp7N7TUNAJxFQGcmV
7f1CSzUP+PGloieHMqyPeXDbkUhh5eK7zEaufS1HN29RuF2RAylrDdcPwbxW5jkO6Wly0iLlQcZA
jDSpJC47opuPsY7KepESefFg2gFLmYb4SQ3EgiDf+aOZcbbWNFe6IUrU4RqAEOMjLo84pozZQ45V
yUpRw7L69hhzYZUXHXqOqwEN7eMa1IMLRDh2D1OIIviNqsQOqfjsl7qXBB2aCX2zXBCDqkn/v0kg
MMXQ5kqEkdb46LwudOfOcixhkATkHDw8ydaCKyQSMhhDiq+3cDofNkObRB7WWIZq8XPP4eie7ptS
rinfwr+icQ4yzsKe9yPwx94VgxYoFlLJCOE6XeCMN/g8avy1TPSKcVVRyLJOn2G/dQC1xuzbb1Gb
dlxaKZw6uRrrkDYykSYCqdA8j25+Oc/PcVzhupUYv+YZQYRdMZkknj0EfDjMKoyXvInap78Dlyid
RFgKbQYPHSxJX/8gJHkuKWW1CrY6iobRDbTLp1XvYVER+mxBI2kEKGPKwcZ9bOkE9DypSed5fXlq
plK/jFRTSMtFgAcp2/4csRrMfC7/EUeVsSx/Nb27LiCDWQBIGPzANDBFMHSPOx/zXtQLMOV0g/2g
GanytkJLSSof/wBBtVo6JuDqua1QDirqmPcGX85ppYU+impH1QPQiZyaTNiy8yp9O9gfAYLUHvWj
oMeq8DZ8cR3jGtpS1D+alVBMsoqlohLQN5kwGWIOwFHnApO9Jz3WgIMmdjrYVFF22ach/v8SoC2J
ByIdh+bSislv1KdYu324iyNv/9RQMI9PlWnHttej/DF4P9ZYZtuYUjvC67bQW+WJTvHIPgtWou3x
5kGjIXTQJ3CQkErfBHTXck1VSl54EaakCWBn0J45WMTsxX4NgDN2gXtp48oGv7c7mgdU5za15m5W
gVmrS7v8lpiOi9e3DErNqf79Dsq+AeFeHw/H3f9EgnoS9+9Cda8ObGFENxwzu6NjlFsA0vcyo3Mt
PShtXRuDesDGU4xLUPS4vLTy/61orLPZMDuUntzz7jNaX2iO70CCnR0PF6krwHQf0aD6l+sbbWmZ
vkJNUwlsWyXA4M3Eb/kkEaCWom3qe92BJpAmeRmPfjY882oLWeCC3d8ChrvxHnzGvtdg1rUOxb+a
eTSWCONLn6BDJkwYSWkNZUwMxwS4Ih5vRjWE0K5kKCml4YDXagEb0kk/xaXWyQ1POrNq8Zj1rbxW
zbcZSelm87JTGaBwJKtxEWMoCHCdSLJxoFD0It8EgMekk3mTlmvdxdig/oGAGTz/0diOWopB4D27
m4zw9hNxkpleEnHghXkreZSWIOMx6+0bSqukiXNz0yG5B640ERZJCZF1BQR+LbiN//feXkJsoVHq
ZgcgBE5haFvEpSCQu9BY2+lxqQ31cTSVQjMYis7YJ1/i+GMTzVq2pG/Fh9NO868/jT2yVbTOmEtb
+O9DEPp7hm0HVFWLbEfXNsoSuEEM2n0HeGiZnoVGymfnWPoxonDU8IjLv+7qR+uaoBMrLnVrNs7Z
arR8hCsGuoFEyxlDYUaQfa5u+ES596t6/kpTLZazKHUy5kmoS7VQPZH5gNT7bj/k85kyvyraMgYe
zX5GZsxJJdbZgEY/6rEE5J2SKOWrGnuJFx0A0StfkOX4K2vy4w7YrLf8Z3MfBcA15T8gb7nl7PIP
/uhFXEcl0dMxlcneOn6TNdaDRH7Z2247vlDVwWbkxaKh5aVZjD8ktwKEmyfAHSXmpz7hCb2CR4sR
RloQYKdHwI4/R2KknHPmuDq/uhIlVY/y5VqRU5jJx4Zps4KppMfoQwOzfrhAw4/KUB78ym8hKwsU
W61lNbi/cl8+pbpji+VTpQVoEm5VkhaS5TC6VvdSIrPJNWm+S4D4fe0WkMiZIuZ/Np0G+2r5MhZj
4uA2daAZXWSrGjr+Tacg6OlJj/kMA56xpVOzWUAcJlcW06zFchRsKHc7yBRZn7kIepZhXhx/A4uO
OCHqonElCC+UCtuQWuIbhzLIzak/e2mRHvfyRUl231XKsp5D7gPmyFnjFIZNg404DWt9DqtIVEC8
0K22+d69bFZ7CTk6BXO5/ZF7xZd38eDBUnCRegHK2vZaDARFBnDEwhp4pAst5IzMxCGbn1ikwnvB
+i9YsvriCTk+s2v6RHm3MRSAFaP/u2HL70vIo6jEj6JBgTYbO4Btk8vK8egAfNudmZc4x8H3ADnw
mT5BIMr5J2cdNEnaAsUcmzgerjxaFR4R8xX/yLEFBbU9aSW7w7adKlfFat8r+tWwD/M6M00u7AB5
gSkn2tU860wpimezCXtRfGEaxP+T8ht7IQKF0YwgX9HetP1ZT3V+TXGLIZSlyyYsG9qxdMuP11KS
l9I4YTsSpDQDpsOypiOXaaEscKVKmlw1PIjuPbRLBMEa6Jk5hgY7NC26KRM+9UG8weGGFe8E5ydD
0QkSc3CBMDXfRsLSC+kErYM4rMPVRi3mYHEydCMrHjOPGthgosqni+UOH3HLnIAp3XpT3+6u6MPq
H5HE39LFo9lVdytwz6bes2bdMFJuVWC3fVAb7NljzeZdVgfdihdytSiKUiil6u7AYej7LHnUqoPS
6+9SyN05Gw9od/QzWUUkA9JuKrkUaBVqPs0cgOdhqdVShrqlE01FABTcsOPnyWSpOYklCAsVvN1F
cRB8KZGiRHWquOx/BECF+mGElWcWw7YyD7watbQF4oQRiJGx+WzBzRidbI+MqQxoOIlkX1H5zSrN
MNSu/NvBi196vY2mH9QvEuydmZFb+8HR3WXVkFhwhpz2fD1kmAFrkQZbjD44es/IIUSSYldPZzs6
JPF3CBLbUz0cRv48eTIgWglJD9q/phw49Z3c3KrtX07IgnUWgw5mNFT1UNAxeiDUK68H7QG2fZo5
0QFTWcu1mmHmb2zwWRMWxYpeNfp82O6bLQa3XPn7Oazn2elYdC+7AiECpu05nYqYF2ZZG4VPYleb
Of/RWLah6uzeOwdE1wwoKApsCS9qjCpFSt01hYD7ZuXVJY/VTw67n0077y66H1727e8dePojmmMr
1rL/YvcT7a+jqwzcsrYOaaOSk/cxTrj+s97PB9YMTrMz63hZgiVVtUMhxVK46o8YkoHIg0AgAg3f
1e1zLGlI1cwFxWQRuM5xXsCm4It1NOqPM4UwBETQNDTbX3KR+CdclS3qL9OycdQcK77K3ax/0ETQ
Gnebnv09jSgiJ5+tpK/RBsic1UhFCmY5JMJOIBPD8y8en0SSbcF9Z55aYA+bhEOj2BPtWItY+03U
zkXhKLH+rw08KrRjvkizH6yvDmw7he4hpak2zdg74kH2yfNIOdV9soL0waafcwsLuN2a7ELNybhx
un/c6MZ/oTpUJmbE4RT01qZhCGBlkdXWUSNfWPNrizmenNb6ZnDFsVaA6LTGyxOyPjHTmo0x6sUM
Iw0wFcWPlgrJv2Gcap0qXz/fRdVowIPV9boaVON08iqG1sihh9PKaxw9RTUCDWvKyDpfLvcQp28/
49s6kgV3APb0rNfTrfEI6/rqpdG6GEZNkaugDSBCCtbvpmrTZGkZ9IQyIwFculDjF6CoImwXBPPa
1KP2y8W8RL7lDGkx/xZz4oobcJ8cLO4z4pm+XnS9vseB4AwpkLbuyOLXiX+RyjmqMFJplPgBPWn+
uWuZEpUOXkeio0F2SbVsfFN1vShyDdqOOyzY5/o5I+dATBtwp2o4TYim0dsNa+3X5OW5GPNGGWm0
qOto9F+dioV3u/aqGlM6X4obexgEf9IGbTXleprOQ6mHAJTYDZ+8T4kciVZmZCd1n8xzaLOyrqZN
NJJDwTylmG5Gh3AfzeGfsj9VZ/YvGnYQlqgmxcZJNpVHndaWUJZfUvK4ErCKQ/6ft67bAKDL1P9P
+tKW9aSn5pZfFmtBANvegrItVirwhNVSVh+xpk8TpFM6LaIjxAc+XuPwxFK734S6AFh+eA/1C7uv
mwgxTxhZ6Yw2T2HC1Q/8zUt8Uw/9mfqYNuMwvkBHl++Jc/7DHETs1jS73iQFut+YQSXCRS1cb3xt
YCKE2412Z/QBKjybUCbOw7XzZQxmAhJNfJDFH3xwfigOUQ2sBTFtCNgpxzUuiC4W8817PX3HwHlp
KvnoZss3EEovhIjkv2rUopPUSAIyYrT3oOlgBhzOuuIHyqpoI5tR1s/qru/05knnpLGWkTo65jgs
dNaN0Lo5NQ/9vFMTEjLU6Mg7ApkEIqsYWf0v7YipAAKpKmYjLw79wwsr2zR0kx0SNzeTVOKLVPi8
Y9utRNhEj2CZ3dRsbVYx6phkmYtHUFjk6AIeLZznTzgLMKGQixZv6hMCvkomAhojJqDRwEKa713t
EqwydZz/ZAU1m0AS2oCfjJmYkwsY1KlcAFfZQSgD89BYIph04qVW9vitw8fm0d3ke7ToiIvcKwbu
rzP5N1HW+Kw36nzA6oSiiM4ZE3X60xJsEqLHkUl+LXn75ETwLxcFl2qw/S/Z7eajdkyjkosFZdWH
4OCKay0YTVfqjybRceNrgE38Emg06r9qTafY0pDaM/taHrcHX0BaD9Z6zpOlincsXXSNkLOWXbAB
JkP/YjbalcT9tNA+iPxzq9EP3b2piY2HVCK7rz/iZilvp1UOscAF5m1O88skg0MfSvgxXHWVTips
3fTkSW0K/yiOMiJd8RLO3Ii2fPB7riD21W3WpAIeaSTyPxuUmZ5QGCqE1usHWZCJQdOVpgcOKHKy
oxOoILWsV3p6iqucBMCErl956lBNkIqgvn5kh2BSdI5y5gRuYjufmYmJLTeuDuEyvJjN0jneoN3D
GOJGqEK1/Dn2QzHLeLogYvyarDE7kiIH9kdNsO9tVw1voHGjzaYmJ5tgtunIAO77fJIKXrPaN0zk
a8GSZKroLUFrh0WmY4pnGbJWxrzi2QJrCMB2jJU03J7M603ClnpwRaZPKIRAsDZ0VwRZxxbj6Ru/
IbKV1yySJlErDU0IiUb6GoyBPVgZ7t1X8jegGEX6R9HHB3MKkF2Yijgpl8qjnwpGF9H3Nfi6WWt/
cRjK1ekLwHaIOs/+RQ4ya59MmDdtUtyHZaGIHAeS4Gle2CvPJSi6CFcRsFFaCxAqUdieBj0JNfKF
TI0kq8jxInaIAz+xNNTEG+9VAUvIVo5vBZmbOYKfoX6kZ8E7UiWoHVAClqzwU7eJmcGcijeqs9t6
k/hjKHr4IbdsefNPmjuQsdyU3tf7Vg0zFLGGDaZEe7uD9Gq7+BOkEQ7Dne4M9UdtKECGR130gNh6
Wf9b3LbGLNInpxaVk+xwQTKVrS+z8myH6bpSRuP3oM1YFnFA7zTnVvtiFCGy+CF/lLB50nZ7xbek
VB+P/iECBgQN0ePtYF+lRojcftRsgkgHkNnxosE17kAcAWi2RJUfzU33wg8denTAYu0RWPhjTpS2
woeiajupPsHAMpYdYnc3Y3B/gSTdmx1rnk5cxpvPTVTWaJqiGKpjd4DC9pQugROy2V5uhhSZmDJb
LSMX4CJSZviykuJCM3sj5ElYHYJgia2avMK3cDI5ap8jytknM8KQQUY6UlfhVPEpB9XeLCr0hCDB
VRFInd1Sp5O4OtiCcKThhEsds4kx51u+CkOPaoc1UIFsW00tC40VT4z1CK5rHJhiakAPTwPAQrdk
08jJV6f2IpNKmloNiT5dyPA3L+Fs2rCtdSItZqEy3bp0Raio3NNYZdb3wTwOvHRqn5yBDP60jHh2
lEjyMafIjlfZ5CdNPziqhLDxSVnj85+uBB6G5gTj6yZF+gqeN3vICT4Nr68r6/XgJiFY7f3oZjxp
lBhwTohRXpEOj6jHwR7qD03HXRUpF9Zxt2FOoERhBDGZPZLZJ40nYtF8PUQUQPEdMBVZo4sJJXwG
rFnPqrD1RIEEmWnuISWjhspbYJyK/wU+LBoLM9FifHs3ZmI/uJGEedVMUspRp/GuEZSldhhGh4Gx
gvYZqTKcuiokE6VPHP9r88zaPYBitYy7p2F/FOGaqvrV3U8ypjzg/3yXqJN36+wntAo53Ciwyick
f4r5goDJJyGdQKMvlKrkIA9TkCWFD6K+rIqaof/vdRyor6JMjF5+6u5EPlUGwUCO8O9XX+aYW51H
PfZEovN/e/ieMxDqH+lMp+Xp/ceZG+9iU+cK76RTg1nJPQO7SJLgvZCDewAFPpgVueU42jxk9taD
Uzij9GWZcW2Xkc0AGdNWKll3geaQa5vBqpPcfzxKM7WdrNHec//G44sxpHKxxx2hPWd4aO8vdbBO
1wJMHfuWlGO3ZA04Soq9CEDSoieWIMM+yPF6ZbPX4LJVdtnWOUJZMLZKxoN/WQhlvVWz5axrvEso
oWwA4yHZTipwtb8ViiewsFFduh4F4jPsKGuLf06wjdYVqn4SyONy7H4R1W2BywvL3JEnUFleQ7+v
SwITBqRelTzTD6N58IAvMUyvfrjWxA4nGLje2imETTEt1pRS6YBR54+lu4HWC03MdmOoZE4Qe4Re
fbqgGeV43gXIqkQcZlY7fz1vG3Q7VwdmUXKOTCL+wfR5mI7JUJNCnhmNi/p+VgVebHA/rNZra/9C
1W98b3XSb6RBaIDxq0U7zZ02GX/kExRskAzMUb4aYoGSCweh99RqMz64sB3Sac0z6n3wCm4X4CuX
hHlzSFa+l9VbXqhFQUHl77jsz0B7tRJpuxiilbb1osfXxJJ0BHuE587VDWdSxfWX+PzDZ3kU5+QE
DMw4aUjUB2gSDKkx4psHz17EXhXwI3oQNfed01N0+MFohZokEut2xsJ+qnTlMIToNupzpO7VZ75U
i0riiEjSGj/ig4owbNTkZ2zjaD6WTjp0JCqW25+JaL7mNvFeBArYLUgVZxozRqBuN9Q90fBJ+g9y
9UUw2fBaArRwK2PvTBTmBCtJICPz7sPBw11K7TkZRtE0lqEXgy5B5RPiH21v/ktIjF8+5NA2mrpR
NeeTBa7QEF+5niuMmgChXrG5qjF7D8566V2o26r3H+k3GVuXd7dLIIAbczDkfH4bLSD7HJgpObX8
udFzXV7HB5TaqDkQB4WJElOZXTNnCc6cWffZ268JuHlsTG87gcLtOFpuSKoUIIec1Xo/Lp/beXbq
jcdVxqgNFeMcRmI2To3yT3bTSOAqjqRHpuyVFrzmtEXsb8wr6LcsNaEzDQySqt1cusQG8Av+AF5K
w8gCypwfaLdWE8a2FUvR3wjSJCwRfoE8CE3UAKW74NuQt/vkFU5ygeBCnnYn16Uddb/+BcP4BUH9
Bs8owZSLcyMnZHjJg6/PCApfqPJZ7CmH2bfQvGwCd+t6xG+kJ8u+82enavlkLZ53rgD3jMDHrApV
I4MqnHMbc42hvVqyEGGISKZ9AZdvx7T6FX3Ae7/zdEDt0VvqhA+gz488KXwjBnK4I5eWFtLxYB8/
iizlPTpkgzQ9n2G8B+DSjFJiSlFW5kQCdrZRvXqQqurZZBe9+5+ADGVg76H25uiLB+Zt1zlQRA9B
MY0LBdU20q7QeYtuvkpBv1sj60yMNsXu2XiulusyOWkGSJVdyuQnBShjAObUpmxmulyNVuY2bH5f
KSGL6/F5Ug+6FplBrgWa3V7r+chiTDUq++zkbACH5GElEO3rJdD0rDJSQO/obmJ2LP7pn/EQTc5h
M6QlpeO6La4Rc/aQ4z+gotNvZ2gLLKxm4kg6uOnsOQZ2zmx4OugyOclOyABLHmanQLtDFPgiBz7g
A3yvmd+bN65YrtpCnyDz8jPghO1YN85xaMQVARIICMIFuhg+mUmajQCIY1sDoZi0jcE4gtN3sPvU
1wk3VYnj9uAFOccBoOv1DbMUoqAVrzYDnVjL3yHhrF0E3/6NSRGgfhn3AaCm2apz3wv8zYgKWXAg
St1crR5CupRX0qtFAzoVcZlzTBx+bbb0Pbnjiq1FDE4e3/KR5OIHLGMCnFWN5PUCPIMP7a15rcQ3
R3Hx8mFne1McsnftaPOcHdVB6BBGnwBBerPI96yuNjQWlsJ47fNp/Q9vgWZONObSbPMnrOBpFmzd
GBgRb/JB7UxBVVpiPW2Q64IcD44rvSmV1J7412Oq74PDNNrERwRo4cOlm1RU927Ftz8SFH8oWjZA
aIpHuXbXPbHBo4ll9ZpqIA2leJRQM0ykUUMomEiZjDt05MEmK+T3YjajeWoS3sNse3B2tAERu8pZ
2CVacq3qBMFoatGwSxd5hTy/NuykBGOFsIU+VN4m+Dv4hQ4gR75qCjBcU9Ypj8BPByzp3qMHGqFm
xY2mIpc+ty0jOFXiy5KlKULxXmRE6UgUEN+AedI2FiGai1I7ARGNun+CM8YsyduBsvWzozssGfFQ
yxHu5cAgzTRShobEP8X+2fDsWKHtsogNXTOTUwShkYXXdfkBkc34UQNdvP1FTpK3aG80n9ICZ1ca
uYza391FgDwxLzti4ClcFvCiEJ1q3p/Kud1lAYLWA5stXBJ40i2hT5R9ey7wdBCJ/T8EEOrBsk87
wjZY7wKxVsuxjmSGH/kaNaAxlfFE15xLOoRdc4rfu1nKBRN7d9OoXhsavR/p+N8kNkzb2f8gAypW
fCLy8TMcLt9TSXGtGEKKFAmMo/aLUQMHhZCgjniAnCltvQfpEj1dQ6oWDoke0guXCA/1KODghRw/
IaB1kJf2ZQr491RYRv8RFiITS6ix/aBaqlFh9yKT/PgstZWUfaLxcBHnVlXLmgUFZu0rxMbu8gKU
76NgC2pgQ9pIK33sS9hXf8GbXy+w+/QNMy81iyJVw/CY1cvPZauquNb0JOZ8L0nBo0iVXUMH5oRt
ekni1FhVMncMSVmxdiX2klCz9mgQ6HX9zonuhYtEobxZ92yJzD1HsxZ385fHw/+E2QUEmPoUcr0u
mRsJmiN2NQoIBly17YjEh0hSa7XQQ59RUNMxQjTgWwuDwwWSsnq7jJGdpHbMVBVF+Xj7SY+ZRslM
2AOQOu0eFne6s8e4Xfs/Q9lTQ+6It+L7tkNI44epHQaI65Q1iZAm2ySXFPhtNxc8bc9VEkWXaNek
qkomHqKbDp49Lp2vQJof+f5fNv831yBNJhS7UtbOcUf5WnPKo8Jyrs2+/fcBWUP2a41PJbFtdylw
+CFyHQvuBMiJTeTjch7rD6MOuncaqz5I71TBuCBLMf/lFKU8KTqYdCFh7dIbakkIukRhPt4NmN2R
1aUyom68wwjw72tiDcLLRXH3SFGSyhQXQh5w6ZuAaTl8j2DhSHdDO3NW9dVJdCq77nD9dhaqgRv6
HIaHQniJsnAuI1mtqikY20SmlPaAqSTwj4mOAteN0aKtUapIDNqbfYHSo02jkvcCbcjvIr3z6/9E
Ilnzq3RkFi0bLjO8T9AvkI+aB2dpQe4xZh4oq6KQ+sv1Fe/6lk6E0FjCOYYUuonPseNf13VRGtTB
CWVgxSOzeK7NuSh4f3FoKSZydZxGbJ+NNRv4m6RiFE8EOo0RFmEXdLYv1BMLvSh2tEZfbzCg1Hdo
iKhkX2cf5y2Ws5t3Kt+ruO4du3Zu30GyzDsOrneN+wh+8dF19esjxd8lmOD+H3yBwJ/udJvDD+fn
KRpF0iq6Ie7k3vQt4/U3p3TIBpk2vDNWApQeyqR9A+Dy7fEX0f9rZ3kSS23kFCBS982esjze783a
tkAKXGJPdTDnb3hvl26HDl3+LLrKfVH6kDon3VwkQasZ4Z6pnHTyMyBEFx2GMcYXMG0anVxwHcT6
FOXvDzkY9XJAcnRXeOPJ9/w3V7vlmz3jiWOE12z1LUYtcart3d9qgSn2VNLyFQ7ruUWdB0wvQDv6
JYwn5AHzGG6xxWm7+Mj6Jo+XjpxxVSa63wIwLK2kxxuiAUQsxK0RGLzbyOZ6QSwf2rUX7Te7hM+o
udNAAMH63hn7SGKMjScTjfwslUEbJAzb4qBLRzkeOea8cwsT31ui5Hl/WKB5NAYn0zDEkQDhOlVG
ge45M6WnIJ1nWF83RkL8MuGDXNjpy42cdCnaY6Rn3B6X/Nco9VG2i/xcNTjTW5H4ZIhcgQOuUU9Q
GCqObAbaPisdc+pT62LVk428GZ8oMJu7C589PoDYY68W/RBh0ehTXiqWJCrPBss3Pt6gCS4Yc0p6
3RvmbspJss4BJT9rglFZEKEVPpz+K++ePZdfnYHc6PYwoQw6CeiFRefNLyRG5M52Nva4RrwP2jLY
gI6kvK2Je7B8g7Dxnv+IGCR9B+q1mjw/3gk1L7K3PnsPwIQOo7rzvvQUPI0WuVEpeZCgMiov7zc6
G6Xt7bmF/Rl5o6pHVpZ3POhi+EdmEI1+3OU1BIRVTKGcTF8+c4w+jASj6g9/kz9Gu92YRREVS2ki
VFGEQeYX7lfCZYN5qEKQzsOZN1ZJL1UgyaLKz3981fLt9oX6VOI7P+qPpwgmqlSyx2d2Ww29M3mk
I3U6t3hLIKmctVuFT5A4r0T5DjGvcBjmvodUrvY+ClryQ8veXEmAFXcMi+eJsyqqD3raMqMAaXdI
/Xyb1sVAb3bEZOrKi2GfR9JqZYb/Vq+gl3xRZxNODCUom23EscMK76F48ywPoCJZ10IXju9i0Fxr
fAZkIi/gkfV5rkA7FqoIKdVXWyUZFn+YIMcyVprQUPYI7bvJXP8BttwnLgfgNu9lUBEdwwiQjamc
AE9OUCu+tdf2SO+3++7asE9YvQRaJrPX9YG89Su5bsJLsNWp+wipwoDpLuyAdfo12rXhFpsaRAmN
uM9XRDIXPQHmq1FCBF/2VAn5FeLMhA2bYOvRKInPeHEED/3NpfRz8ddRo3xV5DH36Iyy66yQAACH
YoF/tiwCqSRpA+idXyMfAbRJsfsnYTTBDIY873aTGLaMMSuquUOVh3vftugpdKD+/ttcO68cwpXV
B0y/Lv7qe6egLC/iGSWzOis7DQZjc7iBRjQKAK+qaMYJ06z2VN7MA/MZ6uK/mqalNWbCdQP4Eg4Z
IfeYkNqBYJCGNUk55IVp63zm3qSXxa9m9MSbQ8e1RAfuO1h09VlwCPrZRWgRwuX5juEoCB+9meB1
R9r1mUDwF8r9Bpt4jCFIMrbFiieo6QLLDTNMMcf3fh9JH3VonVrWT3o8NIEnfAabYBfKkP6yV7Lf
xLPx7VwQ7QKYZCudTw1DEiIbo2rOFmHbl/wmYSfZbxeJ4PA2l7FRHxP2DUf2eEDGv9wvDI7COK/K
KLHJuW2Kgu9iWwNfBTAyIOdG5MSyOiZu9sCXvEQhRJsOsHw+Km9eJP7ic+3VqH1kOymRrS77cGle
r5E0DXo12/rVw/DhElcWen4EW/xlG4Ikt3pk4jRxpxl+wbPbDe/nQ1j0B+45kumNdTJC8u2+Ypz8
Jg4SmaQETuM8GQu/tNc4o+eySjI8VUdI4eEp7DvpqqmAUgtW8WtJtSCk1/z4U0c68yEEMZUEmjgj
8vFZaKvblUwOHn7XAbuWO9xPuwzv1dbSOKqJ8dEIrqxFFXDin7B1HQHgv8gytWeoj52MHXnyG34g
ccZlIXI1BiL35E2SmhCqzCF8Oh3X5KfjvTR8QRX42hwR3Pc+Nw5VgFvyX1tm4XRRboBc1GOLEYeV
e4cK1D8UOFuEFnFEmk1iXDIxy89GqzvF9lSTWIuW8adnsajmAIYUgFbqCxTgIdHNg/mJTKLGm29A
UKRFON+z4aApgvctR3A22gnn5nLCKnZChBNRcchObxvkCHUZEhwfdQ2xtlupDiie+6Paqn7x5+tq
rqsYrQzADe7ApYVSb3SydyCZ67LR5d32vPi8gtsxF2dyhnYwhRoWFbqR8/RPboyFSlkFEyIXF7t2
l3pS4qZ3748LQTqrA3Bq3Kc4ji85DLN5BtYS7q/Q6MYnLFYzgax3DtLH09cq2xMA1zrXPCi6z+bV
q2qlGGYP7NBqfiKPIkzonu9UulswUmvrgL8dgVCfKOi+D2k12b6ZsMly3+Zrd65/wYjNbiF7iXFk
hxgVolx/jELSO9kVKucQbHnmhBkKkx7wunKsWIoRcoZNaUApiEjqqSa4n008JdM2rHE9ixM2ogw+
fpzSQdBtODWNHxPOwEiTmt9ADlLim5rt7GY3AXAxk0H37lZ3NZ9vCNjyAUwu7vcSLoW1orojyE6d
58DutJY/8/AqlQ2VWEUDX2bcRBqaU3Nnw1kb+mpVE5TxmyXGYaB6qGUl2caz8HqWl708yriXbkdq
Xc4wBSlAL+WqtPsV5flt9wxA9AdrfoXLmopkFyFqS+1kueaUL5W9atQA+TGqpX+1Neve0ll1HiTm
ULNiyG7bHLVq/vBitDtoZXye4wcM7WBhZ+Og1BON8LOeBQvfQ3ZwAppa93EQntGYz2RHcuJJ25r5
3/JiJmD1S+sJ3FAH3CYmSRYJ600009a3yhqpYZTlfR93gyWpVlsE7Xd92rYUcYqdGFcswsp3NwFq
Ahu43yS3fujzQ9vLlmL9QiFlyhA3XiJ+xu+9hk+s+wAu2fxpl5PAAHN1Avgv/ag0L5hphp6/qj7J
xlelEhEufuWE2obEGCSR3295kE13ihCK06OK9NI1cfm6Lmd9spycxf1GTJCrJi5/F1RBuBNwa9B1
7sCDFrKXMgsVXQdoACHuvjYaonV7tO8MlFOUsiG9zTzPTJKar9ODljn/R1ZJU/EDCd9DA1XYJfh5
R+jqt0QZZMYX2tE46frafsGOEbezhebrR75pVG4JhFjt9Fxdhd/t0habvAaGLZzzmVc9+vmgXJUU
4PVSJlCPal8aIzOfSkvxhS9/010NmHJxSBbxIRTcJz3nMx+rVq0ik2NMf5y9wBV1BRJse8jguTxV
yN/2s2gLhNPKw8kz0sgDTWXigAr6ESMuQPKI4brwhx2kq2Rc4YN6K7GCeVqPaUOcYxiBJtlMaOei
GclkKHCdPfK1sTlRxSnKlTmdQ0q8aI/Qu+Vi2EPT19MbRKaep+8Ati572MrPXQBorildAv/VWjiU
U5L9xAZuetaAgFmNB7etGMypgKjjHeOB4/TMZWrQ6VYdifiSHLDvyG4Gc/sx7cFlRb+NV8z+/FHY
ft0E1KXcfgihn23tZN2eOfV5j6sefJ/5IMJ+JNrL++9RnyA6w7w2LD0cgFcavMTN4muBARZ3H0af
eK4I0M3AkbiJcBghEQ2YIuKSsVlEB6HdB3tq3WRdwDc2L6jdr8KVPfQUZuYLoojbJ/urPE0crmj4
/p8qybno3OZfrxmnlX+bRfLBTq6N9/Z/n7IFYP5Ovy1e6UivWvvNe3JcRgGFcraSq/JPEGBDW4Ho
/cb2xJDOsGp24E1EbLEQnqQZHUSQJub8dFljppzO65kTTXFHX/laGfyeuMctsxYAtZ9AOd24S6rg
8Sw6mGtkg4Vx5UuCpLiXyHlu1OT+mZzrn6R0DNMASHZ2QnwkWTLmjGVQygWaxls4XYmRFN6RnErj
ZEVWqKjJJ2E1MMZjgiLg0HHlPDokVjPbRGeBXItcVs1X1aALB7redZ+2ZaV3A4sro4zkjkTd5MLT
8uL8r/LDRruw4adS4xQ7iYd6PLIGL93y1Z3tCmLhLk/aiD6PEqtIf4p50Vx4xaSDwPcydbYm2a3p
SQMu0bKamrqGNj/sXvIT3fDkewy7dgKPAdP+YvNsOVCILg7fOYHylB4l5kDBLMcn93Kaf8YIgQht
84+SuVrUGNBBDiOfAejQ1K1Tex7gx8Mr2YVLBJ68hJ7acGcazuFVZ5C848OjeiMtp4CCP8GYm6Z/
ThRGgwpoCmv5F7vFzeymewyRt0AKnnpJbvvI44S4o9OV0NLF4mU1OWwcAfa7MpOExFdi436piEnA
inlvU1h4F/NZB9PPV8vPJZHnDFH55lbNcWGjwcxMyK9JjN+68mrH+xkOI/tLPXdEMcEIQFT4jSV8
lc0/m6sRTr8DlZI+5kck9KBku4w4GA/ibr9zEM4MrwMZCwmVruQTzHTfeW40x2sdsG5feG1/iCu9
z+mcHRJOH4TY334BTH9GsvSJkUAJaJLl+0j94fX1l0b2pOxktIqQ0dLU5ygnOZDUHDdRmX3NUeBg
zYcfSzV++Y8HIHxoaIVRALx92HMqjG13BWoxgaR5qMf0O4ND0l3FWJ157bneYUyHWY0Dz3upf4Ix
rksbjhxvadm9F0j/iTAgQ9bdAna2UF6mfMs7nOCqLSu4jtGNIqo9o9XA3UEfVYDTUzA7lQb9DWqc
5CRZQvxW0s/q7qHUQfJN3jJfGK0kcgsupXnAnt1NUS51XxyfFDDkfm4ZpjEwnz0Gh+t3ARYEjFlc
WxfYO8g9ozadt2EAZmw7Y6de072owOAcPa/9ItUrn4N0je1VMPsEJxfW6sJ1u4iQ/EcGtQlp4GfE
V6Kz4NFZAXZR4q3VT1fEYWF+TUWmEcvy+9cutOFD8oBr4hE+YujR35Tz5pDKMBn+JBZUnZsup96V
rcDU6CJdVd63ZmlfjrX/0qgeai/HIHUL+Z9M5Id3whDnnTJTmwUb6LNC3B3P6YmnYTpuyXd0mclJ
Z1qtL5UHycGaZPgkOCosiBdnlyHNuC9scTjWIPFs3LAGDBUwkQKVLzHtr/fLC6iyeKcc2ie/S7ph
yIUn0VGA60wcZfPK1d2H3nRVuPdJgZj2xT/HdVB4bgMc+v7D/tXxdZAzpYzsEXBBG4LX1tQho+Cw
NfGky6EaIKv/uRltzWVKFf8LaS50bIiKWfGfSpYC9dj66C6OpFjdNCxk98WRkYMUfmaU0b1m3KSW
ORjjsJhsTASXhAfXRkX4aepLAuzGPv4Tc1rJyXFL2IYb1U6j9taZXglehp+r9RzeGQoVGOVSEfNP
iszMlz7qrixDsf0XAhJrTfuW6b5EGT9dtY1MQ+AukEonKLcr3DHsKzrluUG4BiSetM65mnS70Fqi
Ylune8V3tvCY1HKYFH/wLhAoCmo3zmjHtdLjW6jjNwkgRGnf+sZoQQmf9UPBa3pXXIVLeACmjLrE
KDQ4h7o2OeCjxN6u7EqnVWCfC3sxPJlg8tftQB1YpHUT6pBpA9vELpVhBdAPPmHNwlh3tMdkZlNe
LW5WT+eK9x29VF4BNCglpG3ZcZX1+S/Sg42izx1d8dMraxBRYCbOA4oJzNIACEK+y+oL+Z0JAbT2
AINwcI0FudUhWW3cuYDJkv0QOol941NBTyW2CfWW0SIuNdjuVt/f03SFlwLzLYD9Em4dy6d64igu
jwPA4nE3vdsKL3AKAcKB2p0Lf06Y26OWKLbWOsJNh3X3LDYaTHjqWkq6OhhUNxFDK8RsyqZdG0RI
2haHIARZ/iNpEXFk1gSH5tNnrEhSh03O6nIDiYFs/BIg2odiUhAdNdaamwaZ3BmNIEraYpyydLug
ON3wodkQhu/xggu/+qYwVROrY4/BdJcVTMOKlUFFZgHbTV535cZEH2ijoPMT6khh4Dewlc4uDFgM
ox1wLFMGpz62hMzax6sfZzEOF6Kf+cPx47LP7nDRqy4nSHT7mU+kFQj2Ab0gNywz8NAiKMS9dBOI
cliPVg7HVuRndhg9uKSEguvzDj9cN2gO1gq1DXLRoybtLsBpUyMMigrdGCZlt/+fOFzeO3MxIVlQ
7CAi6VGyGucI0aGp2yeXGVx2fgKDUkglUIdvs0X+RGIoG74FKKGCAAS+Y6pambXp96vpO+1jy366
bbgT9jETqB0JsANMJ3kzXUS7BGgCk5dYzbesHdIxN5UwPvRDFTVAaNkS1V+CmH5/3U6ye90iYtkC
bVCwj3xiJBkQ7AktW9P2WJJA8oV1dvsBdHXoyB57SaGItWz07zy9ds0jXesIK3AxD4kmlLdmVYwK
WjyDOjbmDJPAcUYBdk1M4nkrTqNk6I3D9ApcvVOhQHhQh3+nT4qwwvnDwOIHGZ/StzV6o3ZvhI+R
/jHXotJkPCpcs33cOSR0WqxLrpN+YifBBCkbEGA6m0kBowHwT5Adm6rNxioSgU0uauLrnIEUgbN/
1qBlg7CnRQv/Z8sm2Ta7iF6VqHylZvfeV1GqAcjHXjTXdNQPZ0/eaBZfWFkKV8yQsQKmcr5zut09
V9/iCINJcwISuuKQyKjXallu+5uLBaJtt3717DSlV2FTSc9yQCxDCKXUbacn24x6l3ObDxQm5WgA
5iB7DysP4a1z6Q3bsFu4TTH9L1+CrQSuxItCGDZDwrX1xev8jloGbBkA42k4tC5yXBBVgSuB0369
dI8U1WmW1yD5avpbHLnoiPszJRJ6k1qIRVbOMm7OsoaTmecvX09GpWMJGEgukghn09xvr54U4x1j
Qg/7awovRIxKdoC7s4ku2+OqqoZ/XwFc4Yv3VCSwBjS8rip8zi/rHJ0+1KFN8Ohp8PcDrEf64lKQ
0NUUJcmdT7XNVZP9RfXOl24n70T1rSCSX0jCv6FvgrBrh6LuNlfLs89yoX8HCoF9mbzeIIEQWLmw
YugRJ8nyowMOBcDBBLz1Ofgzl5CD58B7Xo0Yl5B+kJt2iOcVdDn4Hl6ifT0I+wMGcYL30C8xi6uq
KsWfQdGa5Mw4s71YyTCUG18B9Gm7dn4gWUc8dthPx0by/E67x4nzP1wcbFfcP7yE3DqTZ4Pi0Yeh
aDlLp0UN1lDpqpBwOq+fqsQQ3IQXZ+mo0bbpLD02b3ZnOvgPIgxR21jGikB8OCCoOw0CwnAVfKHj
AVTIZ2H9w8vdZ1C413G22Q12wT21DMR83PLcjJcIMi7MbhuonAJCg3Oh1hysdXcQqeEbE5jzRUjd
7RVjnFSQLjyOcAPh+TIAcT3JpBvH60Yp2k444cTz85LjAYOlQvQEvqCk97s1ItHr1S4u1DngJDPs
xYy7/6CBnggT+ZxBTO/wqs+PNEZhtUMJERoLOKLCfvBEDVr5qcFjLiH55RNxGuXmdk7I421aiVEf
gj41uAXEytcR2RByQ7fP7Rsdu6yk6etFZdF0QeAYJdMG8gJKaY/t6xbtdcYhqEo2D0/Gs98bTFkw
KIsWGqd22AJXuFY6lp1aADiQRvrwb/qiDt5nXYtvkVm1bQBOenTbAugpY3ZuGAoSrtSditt1/WCN
ZMnCwEVhlIGABsqVeKekm29ZXN8oSyuSZzEuMnry05YNvloOGCmtccJa22A2E1kr/ZG2FLWOTOyJ
lzsFcjIKs4SjUlzfircVvrlPBL8AHExUarCgj6YUjdul07fqNj64HbNLnY3EdW1RWouFX4Zwqjj5
U5HlL4WHJvQjuhpxbdrlYIORXDoNi8/Zn3YA2uJkIvfadiCzum0pFvZF65Sm0lPDPBLjYaMb7724
8nFiEEdGXQaaYz6tkmk8mmHAv2ytEtNa7cmeykx3a1RfaLYwM1bWSpSPvSEiqUFOMXl9CSrNIrSh
r+gJX7d5kNgoz+wj1mXhPLgLjj6HabKTUdKf9eM3UhgeEIRl0LGTRDk7PzF2Uf1ifcmflD0KTYJ/
m3OTCpkiRDfpYV7ZpqBMJASZtvvzSAH2bD6xYZcJ+F6LwLw2R66z093ezX5MwrBhECuQi4UyKI8a
OK3DI0jC+1PnpU7CMunXuvVTNzQOJXWqlIeU8xysl02XLsPUWS+rl7tXG7NtqK2BqDkkYP6yHHu3
T4VzGpLXTcbrhBQxn0OYjbScAhJN7ByI5ptcRQOiR+NZ/jynMzFO+piiPyTV6Uk5ejPb8ADvSRxZ
ojRW87FZlLPcMUfNbjSQeNn2bUxjkejf9brPXSPlctFeY1lk51RH34MZgZStqMGgdQlhZJ8J/9t6
esXxjkIUVImJWRt+l1WWtvXJLHR0qp9PypTYZW+jwrUvftVG1orhQ7p9PczRXQQBADgGZx37b0Kb
fjA3bbwDDO5jKoJ97XY2Pw185nZQYtathM+gyLdJI3kqZGsgrJURnRn1L8WvANrpJXUPO+v42j1a
Fsvf41xXJNlwwfoORBOalcfQTo9EPmmSbHBIO9quvRO86s1mv/6vwx69CjY6Lcw9gG01kuO9qWJE
Y6XVtaC3Fi9zOc4vzlsfWAKU/hAhTop9PyDo902EZnWzXbTnURhQSa7TIhFZgGas5PZMJrag+ENq
weerT5I4FvPtN9iu0Lx2jK8sfo1vuf+WIBKddbpCMVEEJ3dLMrvwo5oY+7m/AhiaFb70t5ZxiWk5
0L1Bu+Cydmr0kiwkudQSR61Gx7UNVWFsmz+shxJN0yns5z0hmG9Fe/zT2J8oAiXMZa8dbVNBEVGn
ZicZu7WVAZlO9y88gPlLgI+4cIxGQUJFxflT/seNUA7gZO9IFbbTNQiDw7WxOoEKIVF4uQ52QICB
X/5nMksl2/PK0lDRdm9nuRxtIwI6ebeTyTkZj3I6FOrPi/QkuZvtIzGssRN+4pEfALrB0f8tBHPw
sgf8nVdpGTlRVhmqN5T/T1PBgGkg++hxju0LBS3mqFXioLE+g19cAv99DwW0SzT5A0Z9v9TmCakN
zi+pMQNpeJi/rTQdKYpeBryLCIsqpI4kOZdszSG2063lOUExfWaOGJ4Y7dyndA1ZErfHkWGBphPH
8O2bcZ4OBUUeroFJHBr9wfqnowPqp6KBWbM59HGbh63JDv9pPjOKr7NwVgiGUrUV+J85I3a7Lj82
WgBo3/X5OEeN2Fgj6UEsdTFYeWm243+vAwj2NUt7lEdjtqQL71eRqSE+Eq/ZUWu396sGaqhiqiEq
L2fO//qF8gG17bSCzzdjNYI+KQv7X7kpn7S5fi3btppha06jM1jKG5BsztZlB94vZtbBxnQ2asZy
2ZG/OEZ38FkSkCjUx2PC/zY1U0F+5f3hYLot6eJoUKY3OJp1hCjTY5rAcaVyc/I7C5a1dLTRHUTW
tmDX+bwt5ZKFJ2D89PumwhqMho+7BTup62UiQjl12EWLin/fADzY04f9w6h32RrigTJks6KeqH8O
J7GWZ5b/FTFKeSvfKM+SDLUN2EBO1N8cKEsUyoeY61JG4Cr3QM2WI2SfbZj4Wk+m9hSHzDm3kD8/
etHh13VqBKz2rtgdRQ3nPWIdbugTfiJP9kzLnKzRE68sgfCsT1lresZoy3sQQPYa8eMgO7Ja3+mm
y/FuiRyHNKHWjmxu+oifYb9uksjBZSn0j3YNMfOiSG9fb3bdutF+aZf0IJidY2Pe3u6+Brvqwaun
/+nppgewjzTxZhr8kORBRFDLbW4rD6vp17tA/obDMgxMx4QJuLG3qB6b+TUj71DErTGwZwlX/FUc
F4oQf3aUkGcYGZlmH3VHRirZxz1kMhaBwvfN7hU3BySLNQxo0gV3ys6X9HdAhXEAnRsoRVB4XQPB
WePtmO7YrlWpi0GLqnCfd6CrAhK5/dRYsfOmBD6ZgqUX4jrAFuIw82IxKx8Kz2pXohfj9KXTvEur
kjlb6mqiHoRfC7F9Vh7OTu3D0c7ZIpkOj1e+K9soaj65ds1lpGUgwszgQDrDpb8EWTjaAL6CCbOM
lhVRo8GKeAdtw41gHjDbhihy5RIRgQiOERMstAI8Pjbh6OXv+jyK8X9OF5pElXMCF/6dQ8Yjzw7L
dHfbX+SDBK6Fm6+x96DuIp6urFXQsBZTBgMB2+dSvy/OPvCE5YeWrocS1O3wZKc+LHBbles933yF
QOclWFQ2QQJN61gJN1MiUW2rP/LTsW+txSwDkj0bSNhdA9cNoRZ3UCkINg+bppa4IB5+0RkC/+Cz
SK39vXQYOzodVJjy46sMTLSwu5AwMQ+DyqF98dcwgPxx3ObXUpxmkvlDkze1LK7Lzp+1is1ZK52O
ZELSMrkKNvscSLfF8nFwogid/43QXjUAPpifU5F5FgK3O9psKKlogLAxaotlpfrzrgd5UmnySQKJ
yIMo570iZFZATjlQxc2tZa6RWEgwudCYiHVBDQ600+0vuDkem4ShTjRWjo/Lq+ztHpKAi+binMYr
mC4DEI4Qw3zNHagnL/I/kDg/ViLEhNKb/42oA1oQ3Ozwxmm99djmjtZEa4tvyEvii5Z5NZJ4T5CE
BREfwU+ZqCP0hqoKQ1IuFJI+qOmDUe9bU7Z7BZeQwqeLzOX/ocHNyPyis79LYB+gmVw2FLnnPbhr
4ZhtCi3gDQrS1f+9VoaF5rJfKwsVJjTKBpkufwGgagC4taN3bS8wJBcD+BHFNF46pd9e5NSuWHoV
V+I/5dJoNYae5gHVPXS56f+g9u3w90Oz8szJVqbjiPsnJ5D7M4CTGtmX7w9V+X8iOpJr0n+EJSnz
aFMuFvZqUyMeVvWkoo9uFMlsxJ6l/zX1HwWKyU386FeEvBgreYgwWx5+REtVJhWkaY1A7u0qIrxI
Inn6yQQwYu1k13BblgggWF7kpn7KEc1dDEIdl2y+5WjdUnVmM3ZZ8LmPdOQzd/CMRChLniZxycks
GsRBKto01IgwN5HxQKwjnSy9Dtk4kXHnOjyIKDJ4kJLbHQGazhYlrv/QU6jPbgx1sDhT1HCcK8uc
y4Qf4VeGIizpaiZ9gyb33vtmpsL/3bfGWUdnsnGGRpvBugemAZPkbN00RdMguazkp7SLFZFTv2fn
pnTRhJgvwqdtc11Mg7F9uvChaeIrt1SM8HAoxq5IusXv0YZ5bf1QwVA3spZip6QtPfLodenTcnr8
qJZ2fRjfzDoSMDNQuvjboSwDgBrZYYa8PQYtjVlSiQHAGj8nojw/cXbCIh1vG+ggfdIW/C8e3qg6
xFw2hgc8jtebVR5ib9rODDbPt2Tm/J3K6h2NcqvzLRTKl93rNUqsu0QjHDTWhrafmfBm9/7eED0/
DpFNZA4hYSvvaQR+GPneLuXbSBLrmuhrHfwvEA30V8JTtV4XBibv6/kHarIPKImUjRCmkFpoBkEm
ZEg4Gr1QbBZG70jrssY/0H7hrIdARq+PusyVeG0RlAfpJFfJl/PyRHQ4Ga2z9wlOTPzDY/BHOpUs
Xl8ieR931DzD+W7SjzFwyO0NxF3+8b32KlefpQgCVIKwR3/SvCO+78JN/LbdXi641QJD4UjfAFV6
URWEXlGgI1O3+KL4XQHobsvrT3talDmTaNXG0ILkX+JT+u+G+SuKJ8Irn+GUe0WAl5XQoPB6fQ7p
oQDb56WnApuwy5Zig2zXZDlzslCZeqDTCDutc92ChcUjeJp+UiqOciBp69IsAwAoQCxhef+2AOfE
M14yQljmdaLMSEIvWSk5BFpAxcRTgSz1ShZuQjm31CDlDp32+duX/p9GP+1EHeq+WKLZQDn60/40
59atWRdICHOxkghNSyo5cKZzjHggAsSgtPrnPHtFmIR2ihrp0coZBvUJTo2MrhRTfCWOK8tDNBIS
MM5mfDAl9j4eCgit+EDnCPDHr6Rttnxxx6S454ktW9xw4mHVvjKgH/ND+pbHhdj23Y7+0uxW4vYR
RmTpnU2hNCsTfP+dlKGVmf+yjenqBa9HqJgE8KHlC6FPi1s3GB/BArwRH10nyl1eaSOpW7XMkYgZ
Cm2h+v/xzyHCHGnQjaT9uYm21uKYGGSuqJOrmc7rGYfXKw1IswavhclnIAz3Ran9+t9H68u9s4Xu
ugogrQOWSsT1PJjFFNp3BIHpFn+r4Tr3h8OkH37bBUQCBawnRqWhF5+YGqGoXbJAkR/fA4ATshUC
37Js74TLbxZGvWbVIkWlOnilSt3q0vrQ6VFV63p7xtlgxmxrkMyYCiUHI5320yFrAHcVbZCHpuPY
RduhlSV903qhshlQiXNy90XOlYLahJl0d4ryGcp63Xo66FZiZxtkIvjLIYEh87MNECr9RormoQ7B
t1T+oSVqXxNEc2sgiiF/vBvjiJnxrpeIrgAEN6iDTeauaJ4UUaXhFqH+UrShoz7NxanPhZk9nskQ
CwTCiBLwfwbkRCTTrCiOt7PJhZiDn0+swci29iWCT7UbFyMzjbOckE8i8UehgXMMx/tV1PNT5GAq
yJbxQDkODgL0PzGSrzbohHUq9HIMCGoJ7i0T+rNXY35kjFfcbHq1/YE6zBdFhUr5U2sa4XJdOxMB
JgDYjGZvsHGoMQTdxWXXGOLiCmJDypyeoMFe2Lpp64tCQtLmQS/WaaZpfZMuxDdBxi4jGVmoiESw
5KumJHT/BN056+TtGmv077ZVu3SixhTY9fnneERbh7lHLSZaiek0fd+XZp5XDZtVm4HgY5Ea3Zfz
Nv0sOH5TVulCSgjqORCtusXspsBAQgUb9dAs8v3fgWNoJ5CWG6akdJWkd/0SsOqNWNYckii2UXRA
hThIZlaSVS929sbjFsufiYjm2t+J0K+p+7U7CnWMFNqqh0tLNnp/84vVQb/Yp+t5xDc1BUeltxcg
plh015wKyrT2rpAya5rvxSJCA48kWHShZxOuRzp18W4/UhMElfJ+WiZSBACzd86ZrXIr4yyDh5Jy
vXP3t2/Sxacu6YwcqL/TFx4xuWnVFBCsPqmRpA8OuFR5lEXDdRSeVf01JvXK3Vv5c6FqBQ23HoDU
bL3Fv3ANkp5PKIKb1YCUpMcVWIwsxmi342uat9XVY+g6vI1Dsa/BAWKFXwIFVyo+fIXXFvaDeVcM
ww2iooHORYJsdJZxOhRqNSUgW/bY4054IeonHwRQoEzM56+Dqs/V+Z3SjB4TwfVtzBTyJHTPjtpo
HGbnO0W8ZrHa5B7x//36b43ToTmv85PUYRXN6LKFY19yv9lzgf76zOzZz+4s7kYI2uX6oFa3I97u
ovDlQNL2x1RgPFXwtgdomAmAQc/nMtz5U2QcrcdBg/F0XKXtcW23IlaUeBQeezxz9kn3ewT3eZiv
3k973uF100ML1JLD0VA+O5tOEoY+XhsUcnPZrGQ6xY8kWUOnufJ5IPhepgigV8CO6SiYHsrEwaM7
FvlR0GunmlIUFhoR+ZfAWeUqEcg1BIx5hGjZVdC3CNVyHZ5iwg/b3g1TqfGFxqHLUwuCYlJi2kzl
A2QV+GnWOwKXt4q7riGUqzU6hWlKHw7O9jm5YZUC1OkpmKOE/mnWifUaaBv2XmYdUnXjl1Gtimv0
+EjEkPPCK09FBqnSbrNX7y9MWXlEo1+SrAqUZzu5bSLEhvnIAR2qkZJrPf8ltR3z7XXT78srMS2J
MzjACzJ4Z/DKwal27x15M82rvip06l4wr/FhPhOLJlSeRqxNprCdMpw6k4riYzWPUllLZm8PK8Jp
H7p36WQQ3fojqIOS95xinJwMGLUAwNu+AErbdvWRFXSzuSvthpOyQqiWGR3aOh/pk/DopbHuXsKU
EEyT/WOAS2Yz5EmuFGYC2rG7WA/1R9KzPCsYHuVIMeJxYMEKpP2MHG2biJFPYlsTaEHJYMVEgCde
dq+d+wUF3ros1J14plUyD4+wML47VJ6WhwlaoMMcOcuOwGtLUaBLXgIT7ckwJWKpq0n5O3MzAAZ8
Dp2Xs6uR2eJzrl2pC+iIHA7zUnwMopJj5gVFrV56uxFCcUy7iKbfn+DaxJQRB3+IFdoRzV16W5gR
ptv5B+vPkFZ22KT+09h1D8LeU+DzfPiZnFAf/Ftp0Ld1TGhadxa+36Doxw4OyIlqo93BPsR4XzzP
y8mnmg1berPYMNDLdKayuO/aDZVR6mlt8NGlLUTpVRTcN/7S32Lg9VWr/fUEa50syhqtrjjWW0o6
4qe4VtNUY/m5ETgwtzK0QQRV50UV+ydwFVLh8q1MWCkKo0RBwqV9RD0ySltHtWAWRNZsSzHQmmCl
ALfwPiSpuKIunLPacH740rfI6CIp9eBacp8AanmWryl6WDOFm7z2M7JR6ttKA7CF6LGBC+TOe7Te
kc0iDU40Vm1OefESeAcE2PKRNLmLiU1vVMaziOjqzuf6CVl4zSB4uR1YvowUsZSfaTJkREELgDfw
389YDzcjR42s0LlUgBgVPcPHqXvYSyjWrxmighGRbUwV2HW2PJoJkqopF7Wzm+gM9sP90tqFO4z8
+92/POV9y/DWKVvs034UXlfyXVPItrBWDCe41aead0ZR6fQ1MzlmsBMKX5ewfTIFCKLw8iQhJvq1
PK2Jhq+E1UaTflGQvbeEyt/ou/eGabw3iNpM4YgOD2fKkPXhOprHGe9A6qJ1CYlt2q8x5te4ev5e
GhCl8RSsREqITlZRb1d4e9ugvJcvuK3yUdmKqUmYx4kSMqpO0Uz8apvERY3hy/+L8drbDuwkmpTF
5rmtFOTdm/7q/U9U7JA3rNP/r1TDucRNcTuuds4lHvGQW6KBnp8GV06H9O3ZH5HC5cHJSAal7W+k
l1ZdxgV2NzykDuO1HcyzfgxHq7QSZhkgNd9A5aN888H91NDv3+0SUVxGRJEmmAfjIb3WkpIrAHLk
eVgO7AfbZUqiSO5qdyy+afozOPvStCyDxBA4el1rIzi4x0p9sQAxdy9tUkkxrdJ1K+TiqdImYr9L
KmQNdTSgbYE+p1hD94V0Ln8OSWCpowwqYGCe7vXDhb/V4BE+KXfqdHVJiqmJ6VmbyKk2ta8IPGr+
r+hy+5YWYehAMDS1fB5qU3abs9HgmMFkxsm9b0LMLUiSCdxcfjwuAOlbxhZbXLd+iMjMJ+u3rl5U
Tx2PWW0RxbepNqW8A/+UusVcZE9DF8MywHtuOcWFw8opdI2nDs6gbhLNxmasad2dhQFISOOnWNFs
k/udu+DyFDwmOX7KzTa1WRHBdZpxH7+iC448hKaGADo3TPNrvCXbl8+s0NMMnLipMVDq7TMZKWDW
XUAGok3CKA/ZewpimgwxslCHAQkblo3DuRMill1shn2Sd1LCViWuzVwPmXdI3RomaZlVNFYnbR+7
9atOvRG4FvjDIf2GJ0UhYwcMu9I0VOXGEKXIbL4/kGBXoTRLCWeWXY5zXbIqlJAcWRehNHghl6n+
UBPkfSRZuMFueClr3GyFSbhSvJMMKB3hKH6bPdNCXowGejP+O3/YOcGPGUdOXaZYeN93xi0o+kLc
anVtEGRGry7feJEcqZ2qm3hQH8IOXbWB6ppBrFkLoESnwsaIPjsqcYYAu/FjEdXtTZmR/cpAMDLf
L2OI57HyPyZWcUhRQ3tFXimNtBr2ZN976xFXQkh2R67rGnNJwx1SRmz82976os4aj5ipChMT17bB
rIbmRwm+c3NtgqXWLfnNMn8iuI/FPTrXqL9IIJ8vao203x4n+75DW32uP10ICk0jP3YZs8h7O8Tx
fT3JPnpSPkz3Krmu/n1tsKv/z8moz9gCUgwCPkIWQ/mXzLjq+XMZHcOVuvyXbd2G+C1LyquexjrZ
3LrocLpfsHJxQJO95p9kePhq0vHnZhgFPbrPtDgvogXzOi+rePbut1xQOc0+4TjFBgKC8DZScbGZ
8pIv+RteiAlHmxI19X4N6bXU6+IO5JpCcOMqiPlhRBt+9S4einZcldSYla6u0bsa2LCeFWjwxZqk
bUbt1kAjPOuu26DyPS7+jDGROjo4mRlYMN5Assf8wKi5ZWo4qsda4TIrcvf7c1ZLQbL2A8IZopts
yGvX81aKjr0amJ3zwpvTwl7ndRbS6pHWTiNo7bdDaDKjv6uk7rkXBFiNoNMR2gCQ15YQ+EJKTLCr
oO0YG2meP3QKxVyec5CtYL94ifV1Wk2HJJYWBrBl1pe36ngKuHO96Yxduc6cSmEbe6XScAx2VErK
WklmqaiFNcWczMpy43KVTTRo//hMdbTWTr+I92DIAvBpKggnH2hbHOCvRdMGDW/4LObQBs28d4Li
H4TfG3fRq/PB5uUIt0HgAejHSbIpW+gGctOcIjLoaI+AeC2pjUwZ2M8e9mJ3I4HwOUFS8MWuvnIk
7m4CdGrA5FI4ZeQwBwE5w9m29vljE21vU09g/8VqFXnHO4lEGyUVrBBg2/Jjhi4Ux//q5Kmo6/1B
Kj8atMv4bN2sJkkH5thn6b8wKDlQz16mtzp2Q5ViYkJHb+y4oiH2ObHJgoDCtLIKkOdp/wMpOZmm
yaUykv/gj7HwYoTBIRvP1/gPvyaXIwHYAPQrAD7tbrMr2c6XPWVnm5oUc+cVueQ6pT1t6n6wvaR4
kl3MIt40Od/Z3LnrtqxMNqdgbf2O3aUIUVDI3ANjbNWB+zrsqFpabJ74KetUDXGtOB+x02vDiZWn
/F5WheYPcTgMGnKiTCTKlGk1f1mlIwpTlACSRZ1fFoE2z229w1rvuIy5Xw0EvnGvf9JICT9XGlp1
AXYhEyYXGt9PTQ6uh+X1VP9oOtNJZHy54M1mfX5YDT7gMaeThd1XII1SG5x7dHT3tgGAVJeS3jmu
sSVHH1sxx5ZWkJxRIrceTZSeIpjMxiUMQF67zV6gJBR/Rt1vuwqi5m6wfI1iULb3Pg668mUznCKz
zcL8k94kSHbOFhC6LiIUOaWUMxzjK/ZM+L8Eh482bqZy4r77kr4angwnma30u6dAQbXNbx8hucBs
H7OWXLJfM628jm+UYuzmy/GzCAVdmog5J2f6N2EQndh9Tmam3JYybbmpDcMPW3WaCh1jz/dy2gX3
9uUcgHMDG3BxV65sIKw3CcGD7bn1CSEGZv5I0Yi+lx/7vxE4CWUBekFkYKSavTwcPq+X41ZO92lf
F6T/66h8TbjdJMDDhLDB9WYuncB0DC1OZWsuoU4RdGewZFyC8ZUWdAamagTp9O0eo3WZ11jsxa+e
Fuk0eeeRQqQrQNsIAhd9VH+s8JZprLoJHE5kcX1+ojfr2kOvGK82KLOUfad4FMZRv6haINb7lgGz
JU6GMgJUfKaDIrtWhmScZYjTSFgx72xSwsDRQk3Za+CgtSrCB/ws0nNUGVnN+Pe6hRFYQfa7CkF1
34auj4z4GP6WOks27EoUQfxZHtC2h7FuSIen9pp6+ZkpdRrv1WcyXXcr8FwHRlGHqfu6ol53IxyY
D8dM1GWhX/l8NcmhBNVw4R1qbR3gYtWqWsvupza7sbZyKecsouNRCR/Lj3LcWpUg0x6AYO1ra/YE
kTpo/p8c8gMUX1mFy3PYSgQgdO8M2xUNjiMNBHqpXR7fTpyiSzCLZqfXAnKOj8Nwt/dqmmx0LRe/
qV4HjPyOFv/O5U+4S56iMBj6lbbquCit4BX+MFF/OyXT8pj/A0qWsCNGr3aVF3Oh/bsQ0y7J7sFV
xtDaNINk1ihMTN4GnwbjgFcucsMIQiBBIX3nYJlie7iGofQD41Ak16F5fxGYAYHh/f6/3PxgpAms
OnCfevhzpmcbqM3qGS9Ni4GDEjjNNI3un+68Tx1CYCBrYv4B6aAvx3j4xo9eRwk1t/MCAKlG76a3
U6M4flgMpQRgPsTjigfF0xezb0J8ZgVfqDlYC2oTHZ8tR2S9aqpY5MQ9kU/2eusdyy15/7ph5a3v
An/HKDfun0mB18oZChwiU2i8itKzoIiMO6zDyDuhvZKGpTcsQQmFQ0/PKusRx1Zx/HB+mjqhczp+
+9ZXsM90VKms7OqBDdJUkhTR4IVPtUtaNQhk5ogTsqvRghLY0uU5yACnHUjtNu6/AKBN5eam3hHX
ILXUAiwp5HLxoSJafLtCIHsYHyMOLYNdxctC6XXsKdRLTZjxSyY/byTWEUIr662ra1GzNyJez9Vd
Cgd3zqpWmf/Y4o6H40qzjyP8Nj6M3e/gkOGSFVxoTfa+KAML1UAOTXJF5uOzISzwAOFHcBt81jce
MGrYQukTYvnfXJUdVpLjyS77CVOH//7mAl8SiEQWX6K8wuKyxx83m9xfQdev5gtdIodRyY4cHK6M
wqDtl0RrpB6bpHPqRVMuBbrgnDM5Ptu9p1CouwrqVdNTMbuIPyM4fCWCSftPyto7TRyNkTiGavM3
oiPkZW01mNmV2vPLc1taX1n7qr1QKSLyf7p9wLzLWRuI1F6vZeR0B/7ZEZM2ibwT4ubONO6qgL9v
QmIj8/6K084qCsrn0byCVnXtqBqrmZCPXqv5EakHwSfglmfVbdVOOmu2HfDbsL9SPI6xM167BV8t
t8WMqUYYXlMnHHjl+0C9p2PFAXCtjWM+Q8jwTek9g0/c8u/7u0O+Q2yfIMrEy9KAl7uCqwDZHkKl
YkQyRA78lq22UzdG3jdhjlMziMosoW5G32xpfC3WnLh1QZ2yY0Y6xY6UrU9kmawGx76nuOqhG8EX
lxQ0NLxToP9ZAGHP6vsN8lBJzb/+2GnC7PBFmq43d9SniHSb5Cvb27eN8jbsPomKdKRewuNCPcIC
Bw8NgZaKT+ylOH4pNE0TzXrubCKHQ2PrY9zKGBFmlokeUQvVgbS/kC9OeNMW0LsJbvG0ycn5ahpM
fii0ufVR6ZXWuyZbGWNJyUoYiGOCx31sBtD2G+z/bVD3YNkw40dBkGPXKni+Pzp9/SuDCVd7Bg2H
B5A27h2gyAFaZNc7sni2w+4wnfe38p02UWTO4kqYozIMrxDBbz9WRGzi6Tbiwfn53GofcLqt/52s
5Z7e+NAxWFew7A1l+k6do26lwyYUccEQnCn7+PQl96L7LF3rRvM/KOBH3vuECpPTkKY2urU+qJhk
a4jE6Pr8OqCxzzzkmgWrI3FNo1W1Q3Cj2T4CHc5jobSHaODu6jkbcNPgp6EStX6ruXxI1ze+ERSv
EgrIBuknE2w2iz/M1xm3dtgv9Eu9J6JPucqDH9DgdkWWWexGtPkmsB1guX+G6XlFzvYzhMnzlqCz
37R5n7+QpDogx0S41K0rXfSTd8Dq6wDUBed9256BCcQbC5rNQAu3BQpMRJq9TMcah/yb3Rjwtrl8
8opTUNLCYo+T21m3WFCoY163kXfq29STWbmU/sWepwjoDvfka0x5prI2sUDROZTTxrS7UGH06WkL
oWIAKfkg6Tq2pZ3vAoXnMh232yFHnD9rtzLEj/BSq32qkDphu81PAyQ0BbBdtci+mx2SUgBkFcuv
JvpfPXt6FKwlpka5LwuGpwfHiXBaFmzpK9oG+QdsCX3jTjh0hpIEvYE8Bdjq90gvXpKvCA6r9/Jn
VusLAG4K3XwR9bajyMCsQXXNsfouUbyZo4j37gB6ROXMDluO4BzNWOJuTa3QBNdl1Et4GgTejK0f
5MM0WsXdS+O4yDRFzuogZLrq/JzW2DkV8bA9qHlMh9jlEu4veyoJcM//g+Sgu+BmoMVwc0hkiZhE
QCsZvN0FmR+9DKBWP8hzEVFY9LNe/rcW7KX00Z6eCKaQVeGulooGjRtVMTvGpLVj+0O2PIDHFxSy
uqn4rHIg7jrsPLGRaiUehz91EZoNzV6EUXa/whDs01drRG/XlNanFqStw7dviABgWurWCLNF/T4G
BFnj+txvLvfZ3EfMwO8aIfBfV00ChHMR7bSJKlUHDWsnoMNG6hKlYj/6L30cZsOr73icyybFZuyZ
rSZAJxqUPHbms/5qJDBVW9HXkPiAVhlHjKtAOwTTpW26JqRlHjTBFc8SNv8HAuqqK4ai7vyw7/lX
nUC2rkond4K7wSlrPAE/U+HMx4hIqCylNwrcN62U434Sa3ltAnIz0Mnfuo9elH9cbMo6tK9Q13b7
Wqu3btS3F2ZjSM8tregKHmWW+nEb9FKvL+lD7jqiftDv+jdLTXIz0cibSpLLXeFJeatDGNegSCMf
ZpSwmdvJAJUjltwCGit56btfb/d8BSuMzIt2NefTtbTaF+cytvD3fz6BRwuT+At6chdTJJQYA/IX
BKhSBwtLNwoFygsmKwVQj9TAaA9GOhknvmJLZKo3Gtm36NaQPG5v3cHkqbUvva8ZNAXBi6w1WB5z
MSBEIAi0yZqeuqcll4EsWsszHigbbonjiTPvvPEyb6rtE/qKXE+lumlKjBOy8JxG4yqKyhOyyJhz
AKDaiWkNtStjpKUI7rCFTaVBeYysLpr5zlayXTjfnN6t/VynCsyUl9qp5jpAIC2H87ICi8L/sfIb
CzQsH/bPNqGFZbCsQ5wIQJkI0V5Lm2W0+X0VI9po8kD9yFaWQno14g79KepCmSbrm3vB5RCHev/N
Mri1ZIxYqRytOUB9uRTSqr3wpnH6qZJcoXgmCducIrd8jLZqaFqryGcVKJy9ztQXGYqnVzNNiH6c
ElNoB/ssibTI853E1Gezw1H9BOFg6NGArFW5YRgjhuQDzoJSAdg4mkhGEuKJzwHcOFRzofu0kUAq
znnyQhrUbpef4l2UiC52TdMb0zm3XaQ3j9kLKuedcCduMaEdsPr4nmjcDCoWwDHjKTaWQPv5py3F
RURJW/fAL2G3sqXSpm2en2WmWk5DnumfhJuBmgpzrzs9CTIjjTg/gqhVaSfMkArnrfZms34n2j2H
tVJ7vjsPd88uYdFj/jrIXCOT8oZmFPS4nlbwK6aWkhNFDQv6ONP8pcCtxFgagJzkRk7ScvkybfV+
vNLkQtKmHJmIiN867BEXiLyMBEJFSPN5C9SwuMVlEKAXasTV20fLu+LSWrn1ptpJPtupj/ThBd+u
dvPozRHx/IcWgY2IgVtutsau0N98EI4/5Xq1V4bMEJ5WvcT8MtwEL7gF0zb42qHCdPzia4fiKmVr
3e3QZYLF/aLh+bYUnYDrEadcVysCHasXKPnf6fd8fIr6oUpHYp3e+LNGtvqipux1P38+zrsFfeBp
xdqiudYfVAwPhcJ3rkiCVwJ+Frf3++6QgapVPSSzKIJEv7XWGCj6mWAuMX66icpSdaQl2cTtMYIh
NBWgmcpgUUGKRn2tkjz2zKnckYQ3e6KdxsmDDJGahtPsWZYz7dMQS94E42qf13fGSGz/OYBTMOnZ
bf7zswy0+dFR7BoDjo9Y5pKv318A/RrfluvzTuOyp53B+WD+3fLgkypQVtdhsyUIqwZTPvK9WDAs
cdseYWikXdeck9ZuJLgXb6ErcJPM4JA0+IlNOlgBKIqJFCy7aoVJPSBDGY562rH5OK1vdvK7Qls0
1hqXD29+4v7BUVUSfzUksBZg+VNO9uJopmkdAXoAql+joNnYQIHvCir2tXhbci+KKbU4Url15DxV
zXO8CmROtkO5c985R8qPLYg4dY6nBb18EtROl7MU89qLVijc92CHWkruGbbR7Zd4cQKW+O0a0KjW
tcSGwi1FTSGKdA1gGXLbvfRwmYsIx8Sb/QxAd6Def0ZFHUyrevWjhkqWp7b5bfe4Imr1tvyCPMpP
F3bj3/qTvhS6Vv3c/xNqn+iGnInFa1ukov1YkUrdhixgecGQQGP99DYfZdXT2PcTlbJcWpoMorwe
gPhYL5wDNO7oxX8impZG+KOVk17G2jSsTtlwWBM6s0DyCqcsvkqLwlwoFwjXK7SocKazijgrIRRL
Hk1aWXEW8iuItZ/TCWPD4CZYj8/XkHYBG89vUCkJALJDIkzbsVAQsz8gjHuPNuiSRCJohyablBw5
P9dwP0R9tdt2OA89+5wt7KSeogYaJAc9rk224MA60VhgfwJYE9X1d9lTenrwLMA/lB2K/dlrWj6M
9BScy30nY7B+vNw9GeOGGDEBz3srgaE4gC+AaBZPiQvHNMqbO4/LI7D9AxdRp5gpXRc3JC7RyqJm
F4qXwe6Csrv4RlemqxqRjjhaYAD9qX+kxhNqTlqkxr9uo4FECeQyVLkpFYgdfHY6PMgNVzb1Ys1i
tcOrnvraYp45DFZrVw8T4K74FUnS3LctcP87DfGGiTZUH8nt63k9URWCe/2Jj3ppvkVoNfTb2FCn
nX1XmphM3o9uber8qctXHNWAR/yLkG6MjMKDInJvFKJ/KR1O4v7yowL9fNKvTg3fPXTlfyQGh3ib
9JqTRimqmqFHNZOgvunDNhdrH30YVGI9v9a0+AGwHOV0TXCe1KrG98f3ZGIHzTmX+zFgesAfa0q1
Fm82xCSf/1axmIiTvmMbqjv2GInIVpRMDmrdxBM4J0UwHtpMW9BAPOCdSD1t6zOn7kp/UKNatjD2
CPUnMeRaVXGTKhV5XaQIesodGRhI3STAIaNeG0lr4s4GXvyT6fxO3cLvoo4RMNdvvkzAoKAZ7f86
sCrmdKX2nmOgX07oaJhyDn2RlcOXNF3262mPj2QvDe1KMXOT2lf9w0Zo9RvKHwR1SaTEK99SvGPp
OPPY8buI16SJFyaOlXYLFG+vQUlTA2LMze5nt6Ufd4HJ0+xiHK20ymecsqmlWqmuxL0OISxRA2rO
tPXtvxPdjuaKbIJsP9fa3MJjjd5mfl0QRCcN4esBm0BJKAjdFaLxCEvVSOTGKUQoRUu2Hf34g47s
PQtQmFyL6jncDuJfluM+vJC+hq3pnIdTPaVWoUSrFHfyTvPOAeEKRoRVrunPlsesRpfu0CVBIYzl
9c7bOD/yGSVzKdrd6MboquphD4BsgZZWCSRFvYSBJxOrMIGri1D3ddib9RXpqm6weNfcOWxmOwB/
+J9eKu9UbAXVgIZheBjWQ/kvaoI5fPHque9rQaUYtPFDG1RKjBSxVm2NpXer6zWm8yYe3u47mKAw
hqRUoXVsUKPin+gS/KEZ/jfZmlRdbzOFAOXIqRlD7776gw1Sm6SLXc/QWVqOY79ZEx0hLAgW82g7
y11fAFQnO620/wI6O482qi7Fmqnk6C/bGkgHvvFOPdoNm4gp2+mwy/mmKbOH0Opl5RT0oKBo88aZ
/rn5pUJFxnuxmH0ipERj9s1J0G/RAz/OAUo+F1RlOyjwLwL2m+9Lk3TxL9niUZh2a0QHZPdhlf7+
+VcqIkgoi3q3tTt9gCUL0CyjLTKGHcJwUTZIJa3K0Bmo1MFeYFn75NhP/cUuHRkb6G/gnmMhVz/i
bhcFU4njrftFh9D68w13MAa7ES7NCURKLbnyLivYIAsBxvvJnKyK6a/f9DbH2hGEY7JoVLzF2XI0
9g7LYLzVTa9aJlZtcPK3yQTg9yW2ytlEWmSbJIDhc4ijFCGyGb61k2We4/fmK5gxgho+Q5fi9jyT
KjXL1Qf4973qKp5rzLHYzzPKg202PVi0+Xr3+WDn9ewGbRqA0K5kY+wByKt1leUd9IhdBPHkChVe
XL32d6DX7NUgybCXZt6/kFk6C5+i3Xx28hS31ujOVghJtzeKMSuLNsMBEg+0tS1lbzF+h9lw+V/s
nx24MkNCZvH6XtaDuDXiayzA7O0/4KHKJXUmHHS5t3uEH5Xy0rVHxq/5D+sZdxpfrE/m+DEAYBs2
KKKkUMa2y1EIaDEfz9QF8oF5LU2j40rKNWpgVlRFPg5Z4E2eJeJvlXwVpf9jNurcCIVefR+KfgpZ
z9SHfwHq2FM1c/Z/JU4NcyPNLJvGNDplVB12WbYWciEanq/co6ZjnXyFWxIfPnVIT1JA6Fj70Fiu
i355nRwhI7uUhG/6SxhERRWyNjljBJQSejlR1F4gdq5BE+eVwoFaMSFopd2rFJaSA7A1QevOpVxX
b9DAMBlSPgS8QY3xKbP7XdW5Xd8SZbCpm1NdTjFf2Yqg8lwtLTxWgqcLHdLaYwHa3V1pLITt3KBE
s/Xsb8ZFB4/tm4tD4Kfw6Jp681Z6sZKv1P8OwOSX3JbK0VYIAG6ETKlpi3I/J/gM2sUJliZ0yMkE
pgJg5XUtyRz2sd8e7cZoGQ1/9Q+c1W63RODzKAcfI9/dMIo5ktVmFxZiCwhAlOx1YeYpuKY4v07/
PPJFL+cViCoC1H5MiO8E6U+bBClGRYBbhDMdX6ypVNvm9hUg0aXW8AoFXgnnlK68dheZyjbbuYhY
s2yyYDooWCCt+aenqDcmeaZ0QK1KKIGds6+1RXEUGvKuW0ykVQgXRcWSJvCaQuTqiFQmPZ7IKIWB
lVEijVLPv6mDvSTDBZquufnNk/UWLuszPM7Xizr+1pN3vbV5aPFX22Is5newo8WuKRVLwMllbLNe
FmsOikg/702Gp0x/bzULgWxsCULpP1UQ/Oe1akpxnQtBhz3z+RUXlZBsldBUpG9nSjB0oQVYb9Rf
8stI9buKUTJC9tOZiQ/YUredEc1ZtnzusWuJkAqMZ2ATh82Hm2B3KzqnRJODUz0nNcJfrOB816uE
WMATfVTlk50KxOxc6oCS+K4XaHAfbYUXyp9AHIEScLR3ELV02l/fLv7JTcNSDgJMqL1VrWystB/F
bPEPWIMGHrdATgCQUICrMURkuJvh9qL/ISsa/OLfXI9I0n9u0Xi1fJkHebwcoLLDZVbbuuCiLVN3
Z4bk5FKeIJsDeuwtSO7S9HvprjooNd99AlEv8QjWiSRa/kPBfgkLjb6it5HNShPCPftc5ifa4Z24
IEzuGbuSA/QUDugvECLf75SBXlb3Cdr7++noHfkl6R17TGIKHlU67ojkCYfM37vi5PLtkbOhtRuK
oDfd6RAP/8HW6kYcujaOmAWP/XLwVU2w894f2TvdpGsT+XkpcEK4QJynTqU0/fMgnXL/N4i1VL1b
5XZ34TuTgxpFkHhvsLT5dsxDHmHX/ciwQTwdNSiI0+dx7DwSYKrxVcGxLxli50RmQqIZHm6hhMnu
YJCqWB2wnb/sFUFxTfMhGzoLOgeCdqNbRhzZxNY8X7m+dYeXJ1PySRoWBCRyYqb1crM43d3YDptM
YhAuesgGGQIxH1qKghA2y/zTrNDWzdYoVF6P4RGzdr/jLq32XnOgn/0fAajIHrTtiGJYxHeCc0tP
Tgj7kaMIB1FtYeJZCqLqBLHiScgwEjf0WjfyDqkBA0ITkNsbwQlS7Vh75yE0ZMnsXSciWnVpCBOV
hIyt4K6GgEOOWUrmvBi8US8FECtuXD0CmBXqgKWAVQ6TalkujiTq/uWSmVCqJABMTMmR9HVshert
KbDwSnVOWJQTNPQVEMfmx7BScKxJLhlpffRv8YlclWKn9rHgTBWN+RNFQkDIyD2fJiNOXavfKo7v
JJciAoMJaa13PbXfNiXxQ9SM2OmpqhbqFA8J3ycmmuLj53PVRb9Bw8n1YilykKa7wfMeQ3TsAu5C
Q/8ARXm/v9FAmqg5z+HiTAIPDBXedNM9ZVOn0posD1jXn/oJHFXdhKzG3Xpi3sJWibPvZ3xPC1VI
YJutyG1lenysorSyiGG6v+3E1ei9lWAmz/5cstL4WXkBeCYl0QqyPb7CodUwfZ5LO6Ein4aM6de0
yWYdrARzMEIAmPlBCu+Ci0YDQBu91D3+JLII3R0oskMOaxuBwnecQqJ1V94VzjhYhE+tRcYNK3Bq
3MjTGwxpesHeUT43XhoPjs4Ui9kNJSlsFExNPGz12mjJzqOAdPA6rzp8pyueI90jEHXrCTu0ipx+
4AfmW0CfbpV2wKhC000949kttjzIksbNreYeTDYxmz/3adfHH3it62t5tMWubbYbSGW0KiwViEpF
Yw1uYJk2LM2EScGYjK4iQ7vq9N4fuSDQA9sHAstNWMEcwOWwh/aimHtEiVRnAu23vY4kH2Uimu8F
FoMYmHO1T1X7Ki/po5rvlv+E0+kNwEHENo/do45BW1uMhfz3jtAl7ATpx2/b8HhOMGIdyajKcwpK
gc/9msLGZk1DWobv2dJALdVsAZMUmxzaqm+rbutjEnfLbyrIkuB9ZlUASiiofacx0NURRK5jJQr5
K+n9g1Dagu58F+i+RkCKNEh/U5GXUYJnFx61+rLqI/1zLAwcQ+jPYgjxp1QofycqmtFpm9gBxL4J
2iRhAfIqpwOmeDfOoamNxTZIMayWII/oIwR6/rOvQl4Y+ZlTohXedn+ceMHYZjYxBil8NCDoodiP
cBa1dX0iuMK03C7fCF3fv+VOTofKpDmf+M4VPxj3guvzNra7ERr3dBgUoRp3U0uoYCzUB5cZ/MIu
dkBD7xALjZGKap2thnfIY4/QhP5nbx48Mp7cqQiwEMMYkBjrlpZzu2oAqL3RLh/rYUghN9XzKj10
DoCvh3KjCvrhXbczqvXN3ziFxmF3drSLfpqr/D7ll3lc/OPNzV0BgBz46uylIm60L260qv7tNI8x
IFu4rWRIL/okz0VEoTQv5ZkTFNFvH2sbABeh3GeVxSgKrGMYYfXmxQKa3C8E968Uaiw3rePzimfM
2sbe6q/vVGt+Mfbq7rDFpowp78hUdNScuAbpCGe2zuaN+nu9eFsSg4/whe26a4WI8SUBA8iob2ou
X9vbMRRp9Vsc52DO/z9/pWyqsrICNWxLN+nW7kcQVrThA6vtBKUqwWEmYy/dtyouRlm4xk7jU3Vy
2ZyDNb8JQcj7NUT515itYYdPp9iFtCWhOKlcO9akoQXm6fGc1R0c4T48Gl1U3vdySZTpF+r1ndAt
L8AIrpzwhQReNktXNy3zsybNNdcZ0auXrNZsgMobbK1ILzMkzrbTQk0tHxlyR7DLe24sx9Z5xuXQ
EhkTtg7cvjKUSADIHdKNecibiVE52IxdMwjkdTG7rP+yWLDBp4HwAxbEUaTFEi3u1/4wU6G7aoTz
CGmcyHgWKxQNkO95IUjXbtr8mssi3IeC/dTHamSyYtxJPR9Wyu/Urwga7jV8cXTOdYoyOi7Bt2sN
fuGjFeSyNbC0ZsJCSeSak7Ie9QP8T8RG8ZKj8inyiBXlxwl6Apg3glpoFgVi6teVdlYgtSVV2oAV
2AQQ79zcVuB3MQHe/8vvjEKFrBb8L+pwnD7NG7gPD/0AGAm54VWRvcuwKUWGYDQImRYmiAgWfXtl
nTciguEdkjA8jkW+IPvfKJ4CUD9h080xNPFBLseqEwh0JFONiI3wKy0JNiUqF1upv+Y4k1CzSB8u
b3CFETZqjGEqOAkZ7r5lcwWkm1L6atU4iUjR0R5Hrlf+AL9V2tUgghVODm2CpoSN4wRUlbzcXd6v
gXXaEOwOIhS6D3iQaOt6Wlndg7fNMUmmaw1hVp8X1XIC/csu3iW36rFux1J8WixSFP+6Cg8cCbtT
kB5m0GeyPl15ncEjagA3+qB+59J8+L0Hn6IB46dwBzk1QkALeCtNCxoBXFy8l7AnUQdaJ0hA8ZsM
hXGhhMjvnNjWkO/BnbMggUNeZMSV2t+Tf8NRY7+34rW2UpPv3xIe3Z0hnRHpGAx5L7jp9yDIJrlX
vV5Py8G+8cwvU8gvXjMKDwb39Jk+uacpvFeopRCwFkkZMICe+QTSfe8z4WkmxvOCrwGYfllHThid
hDyeaVK9EPQ805VPr1ciiBTqAq+3VdI57mip1Mu2KMC5SeRCt96H2V/XiEKz2ba562E5dJtP0QLl
YcrbZlworgBibCXjT1WH4Y9E2lgJtZFo2BPfUN7VXUtrJ3aLeDkvVGeaJVZzk7FBwu1go0+eULYv
thS0m+kaX4kBhPJ+eBtGIaYAz1xhXIl6LQ1IDSYII3UrWIfgyjlj02BdLus1odo6ggcLyC6pgrUs
+Uaa31wu0wZN26lAv8f8wTTYTdF3GZTFvHQMOA2Oo4uKtL8c4olwoYoXa8haEthBxwTSUxaWU1+A
DZ1QTW3iiX4JmoYkglVFbb+5J2eZdKu4JUWfWaKVPsGqHHg/yYBi5Z2XyyjalM5d+vHtViIZiV22
qN1KH25zBf/LK/zIfGa5BxCEsWm1fji61ChuxmfElFEBOGG86inbYt+9X6AjfT1M3bQ8YMlyMP7O
T7Z6kPBhKf1t/IHpGzOBXhuh0ImzR0mRboMLTiHAA6VWSFSMGLeYMcVi1zb2xW/reQlg4NPqdn5B
QikLGSBq31zHDpEYLFCeWYYdZ/qrSVO6/6OKOgwI/yq0J6EQgOv/L1knXmkt5hpYTwyqlwlIsNlm
4MKf+BgggOhGdXghbqHAC/r+Ee8UYwBDPvI9QAE4rzk0hxsn5Z/PD7C8mqPQngirQ2HjVTCtim8B
nT1x8dlHatY+nR1OVR2FIazL0SsBcudgaA4xhxNQFxQNrr6Vlg3btlOLMa1ZDiOigwE1/ee7Ot5t
jV+8fJqnkFZoWZkZa3PW/NLNxqLUbp/wTK6MfN6A3Q7OPcaSNTyQb0CTstYOrROPqbsOmrs/K5fU
gQNNZiw2IJyzlEtzipAtSjEFsc48aa5u1rU1VX1bLrQZsr/bJqTYWTsNxwdOEdLf0uuOv4tq7LYs
zSWz3JDDG8X9NBjwYRboJJMFI9t9fn74z4HAW4zpofov7LSDD9tcFhP+J0SI66aqPCwKKi9fUhWW
c6OfcEvt3hi9KMGZlt6T/9N0GN55Aij1bQ14ysLrhAZdI6lNdmNUUrfPkPEFooFgK70ugkUb0O28
Olxn4RJGvIsRbVrUc6W5AswugIdht9oOORpj5B/X5zbnQfPQAZajh5isO3rrWfc6B2tES+78L752
ILn3waEJ30jvyxTzZIw2BFQ2hPQWvAX7gSbkM4dd4unGqTcyb+k8Gc31JYd1RCi/4rdiVpi2cGXL
i+X70cZECTGMbfwzslGF789jLTwADnV+ijp7eI/lZnXcbFBglxVucsaLWPv799rwuv5g3LCaT4hO
yW8SMCpm6B9kjobE47FRg1dICMyAtqURD8HxevV7D+9j3EU4+B27UjwUg7ck2a1k8DhaZ42e+feR
OP5AgGmXrJxGTYOyWlbb5IKcq8y+tMm7ssiQ05SwravmP17MdqrUndwQOPuDrpBzo/7xB1YQXF6n
Uvb/wO6pbwKVBo/Dr6h2Q/mqYkkAUuW0we6gFC2JLSZqQhPRot+T0hdTxI42X0lb9qYvJ01CxuDp
zZczXmmafF9ecaKKGxIwcOIHOFYd9bJPbYVyQE7qsw+VEjHOz8XY5gVOnncWab6VAzJatWcG4Mfj
4TIj/s3GlgDKgu3wftLlwy1Nt5c6d9+bvjDMC9u0Aje5Md7qBw5p9g22H3NV1P6AtFeuz13Mkn0x
Ad1NIXNQ+Iuzh/+NZ5NY/wDGzPj5VF6GmZHbwQBbIdr6nAVWJCFf1IgCieXuFG1DWQvObaMrBRvp
knWq7K3IvNO13pUG+/RMjz0VJ6nxildgH59HGdjs9i9/Brg904CQhcJtrii7vLsi4IbfvPuCrRho
u6eCoz/IUfBtiajOAfVP70omFb8xnehsUFXUZSQqPvMram5jBHPiexcA6E63rrl1faU1/0ocnbc1
G/AJx6oDK9wCKnq82jf0OWLdAqNZXRxUhpG0dZKv/nIvRKLeUKXun/EJ3poyfdADZEhFfqY8AgPI
AEzdvwi/PN+mspGJLz87mljo/fxcFiq7ll2ERoRNEvXZI/6Byj3pbyY+ZzDVgzI9ZexyZNK/pxaC
M9MfsROyOOiZA9yRkQqgImtiSKpyMJw/3v5Qmx2uInwewTM/TIgntBAn/hcbb74CX+rWal5wTJrm
trKHo1Qj/4tQ/Tp4DMEjUIYL9z+WDr1d+OszcVjAl+HSeYjPuH70PCZzfXclW1BhRsVM5P03R2d/
St5MwBOE3HhcJqtImqjsqUuzPx2QgZIPBgGoV26q/TNVqSMZdOlAXW32CPhoO8Y5tCdqsdu5ykUY
vIOuqqhWO+clPMKzb0tOgNe++0+02OimgyrUnpOacfaOT5BmiR/xLV+N/SuCbGcdKUzwfv6hj868
mKwIXx1egykk8Jyg8WWhUVeF2AatHwQsjE/yiVBLNAyAuMQog8QF9V4pL1Oei+UM6eAuE1SfHwMo
qqSPTopURjgG8aeTZmOe3qtFRafxuPtJ0fHkhBjmGMAdFxJw9wF2Up+yxiiY57AT6lEMWc9VW2p8
oK8JEtIapZrNTVuLkORREEJOd8TRQOKdt+is6tV3Z8PfIde+2OwyofJxUEbISezOpQ8Dba+tDaGP
xZTjRGZQzfATI8HuxQjBQpGl8LVxFymx0XjWmHw3BrAZg5IAZKuZ4gIygxgxsQwfWnPlzsuPv3r6
z+F/OJlYJkb2HMOLlKr21PBlaCKwSkeIuOsFJs9O1vDwLGt9/XBAByGVehGY/sENaz/onnr3sJT0
xHKqkU8fW6cnGry6HZf1R64cEbzHrSk1CsK2BR10wFV9+UbqXSqjiJUBY6DTebnGd0GilxErlNXT
LBwYpylqO/aQKTolYwaDclmpTMLtuDiS1gG8SNywgPYfiFog+stgT26nQF6n60iKIXfSjJjdCwVt
uXu1ZaDLpa/iaysx3t9x3H3IuXduBl/2PWMcX5ZTUhfYamia+kFwuMnbmusY24rN+SzSxIi1Gx8V
9AIvAns1Djq/h8v9TgEo0hAI5dGm0MCAju2dC4sspwPNOnSzSHs7JBWbte8nJExhv2eFOesjmCQW
3+p5Y33hAVtdA7jVE1NHv3pCRvk/dg5BiZr3yUP1rSaVYKcZFGXicbNmZKv5i502rCwGBL/54IG4
loxPt0Cnd112wvOVYohWknx6iutIMdP5/vcZpRf+O05O45qOGbvv1ov4f1ky+eBtLYyKUDaGEKvE
BoAOVO5KOlbj8X00SbynDLGCCixyD5O2T3jugZZ6STiT7D8Ngk938Duzv+u751yhBSlV2D3SBMcs
OqNCh7PkItUa8qsn6wA00bL8K2l7ZzOHj1HuB0zH1IBIrqX86lav1BH+7BYFfJl8BaO0OhlazGxa
5xKqE0ZI6N7wW4giIInX3ON7UsMFmR0SLPDAaKdpeFDfTq2Z6TvxSHDbfgLxLDmfw4AD45WdDYCu
sKDEaNSz1FtBj8kGD3vArDN4pB7d77s78tWUkhf8WlVzflQvooMzDBPBWJRFEuu9uyJvsQztViZ9
8NMr/QHA2ffrE7Ii71IIBL43x/cRfmtedaqmdcQHWjMOIE6F3ZQLIZJjDYF/xLT/e1bqO88OAl04
jEdQMC3P5aDgFs0W7+0MEOF9LSJcWGAtLTCrbMvMtpK8cXj9ItNvAyiXWc37aQKf7/eAaWe3og6g
rqjYMKf5svMaOhm0mbgfEfSvs2C3w+plTulDh6eigf2Yk5yiDqiP1vI4+xwSEn7Hbs/NA7/bR9QG
cUt0Vv1Cicqs7JEtErimWRB5ySCS8aHMvuRvIoZ7p2OnWgYgZPTJx0pjSLVX17JeaFlQA7XtD7Sd
e2W2OodrmDkJnMlKWX61x3REwNEVXTS0UcGxrUZ+GAljRUeOqfqOfdUyn9BAFDzhwCK971hJAvC1
x6WDxRQyDj1NT+/ErtWImzTGouoeqJW0fXf6ZzqEOeIM47mE4T5cBFCBRd/95+XkyGmdTWKHwVE9
CRpvrbsUgiBEukpz16UfNYvewb9/r4weinpPhEhFIFb270HarKuWcLCKyYBoo4UB/pzhmAUmCjsy
snEwTZIRAXkAcs4+YzMjJ4LYOMRv3DAfVBI+MTpsBtIP4HmdboXDEZGUrZUicwos5+nzqj51et/C
ZtJQM9oTD2+0Eec/K7puKvKTyXVsos7DhQ8NEvxBKrVlmXmW6ddmVtV6qEz1jLsCVNnMVhOh5x7l
XMRPwF9IoLHMTr01G+ztMMtwO++m507ql3TBBTfRfAp81CTEtXGtqC3pdCqqN4gmdgZu0ro3aVSy
Fo6GQcHTjJB5/c+ampyzumB45YdwvEBdzg0Z+peqWjxlbsJwwfPfQBlK5Qk6RYgXTnW0YoLV6si1
Bb4L1WvJRsqqVq+5BebkNFtGgufnuRjI0SFY+UzqZ7pPuWHQRwhbYQ3NMdgNGcqOf6lEtCwMt5qS
cTXzloF+GgxFW88IvVVTWYxYhq/HUUARzXA/SBfAUkv0ycPcezFfZMfpVFqyHDGx1uHDaVZjzheW
0nUYiOay7TlmPnlbf0IfNms6yGxPjFuM6qu9Mma9XriX+uos/Tk61xwVjdPrzMrF/6vg9534evIU
rw5tAfWMi2p4DhOP7folu1WYE1tS9kpNY6nzA7oIW5jGQxkoJdw+29JjLvGt4mbKro4fjIXSCfXf
vvaMzl6IPHuFVOC+Szynz7Hx+UnP7Ch8Yi9XyondNPyxYS21ihVeITKs0Fd5n8Px7pCoKxoo2wMY
0Eks72vA0oy98rOGRrUTGg0wsz8Q+xLVi1hoO4fnVBW7KUW2uREDVv2MRiXoYttpBoAdz538SwQL
fVAb+EVIodr1NIeCba6i+NVAX8j8uBXrITD6+/w4eqmIIaXqfgcZpB0c6X6ckotgTJ6bHU9pdASR
1KG/5Sv6SdxfbXThSrfyf8brgH+mzeQwfCx7A5mwcBk45L94VsWtZG3XWRFe3St5s/7mdaixUhKa
hrsPb0JHCF6/3N77mmbXKrY+D+ay40OUjehGgyRmefEPV1qN4I5kjbdBTnzSiks7wXOJnANrwyV5
pWXCrFZgDhgU9eA5iU5JiGsH+u160R26VTkRE/k5/oZIi7o6++OyaPMKoIzxm0LGUxaMRuQpKpdm
4g1WMjLNVBaR54UDBFKjh/vPd821MEEShUtOg8BupGF2HiidFGaCEuOjXsIYq+5CxtJuq9EHyL66
XLI2Tj+lVvkd+1f8h1qFD+PpIkeG98oSnS5JZhdYdiH4bxTwyVt0mq5TDTNBIsMAMzbj5NwRHv6J
ZCwqAohvHPvgb9Jcz/14LitJTTnhK5K6Gn/jAdv0+n1ii/BqqQnl+QKbnhSYPZHPJ56wOOGXdojF
cewPnyd61+uhGIgNdvrtMVGyS4AjtoqWvkjGVwkScNxOVeQWfrFjeSfUwkS2Fij5J7uwIpZ57yP4
7xVpJ5YA/yGz9ipgQP/hvkV6tD5ONCsvS/iMdKP2n6zabrqJRTSt4755xOT+4BRdvTU8g9PACixr
N90KOVDFisD/xefIWUgZ77vR80XDx4ccDSutBXr2brQ9kkdGYwuuvMFQ9J6velQuWC0GvkrY6KK3
+Ii05HEDyGkElg0APZiV33WyBdHuOoTf7rTzpZU4ZJGnKqr9cM+BHcn50HUCFLRWfEaHU6aNwVKS
qFaS8hl+ZtaOJ7WZeztKGfWD4owyvKI8iSbeiX03MdFzV6S+/NJCICw2rNLRa4UhmuWC8AUFn4Q4
10qeF6qmRY7BQvho8/rxrnTblKHbCoSYX+m0mub8zmwbMy40yTZIxfHfsjeaVe9r5y2I/IYxsyiS
P6gpq4vRlOKlijVyxXl5UKXzB0tE02V4+pSPrciMUwCPvUMQy04ssJpHNahDsCrT5uoGPrJ+cLLf
2I6WwghpsXhDXiACQ+dFnJxC38AksiUdLKPXJO1uUEz+ZZr46WcNoHMjaZby3JXmCeDHajIgdxDj
F8QTVQGDtjPBc/fII/hsUY7Lbqyo32G00Yu8qItP9TrFK5o+8sixgWf1pUjQMTil0pRzo2z6C5pO
Zp5/M5zJ0D9Vl6MyNrAt74dg7gpK+htL+9Kdi+jjgHsxnp1CMKQViZyXvmS+L5ZzZwmI/p7g71MS
RXNpgMCE4lmcN78pb1Ft92CvAVozeby3/+SpPBwhqjPOUraV/kMiegeQLPPFFGFx3b3VW5sEwc4x
W6oM1AHPWCzyPAF8F39nkvIss2BjxE80XWJwbEblM5tGd8+vdtc4b8dHmx56JqlfQG0rlQOslRjH
ZGSXA86MCPMUFqZGucxIFrqA3fbNnCrbvZmCa6uhCClNOBVXF4uwPdzzLolgrBDcbGxM/zXCt2IX
NrE9xCi/816AQZ0Qqvyi+6DC/04nwQnbpUKxhCqKO76zatdWhI1qZBw5F8yxwp6biOHPVQuU6+mh
g1AJuD/cGdyyeEaEf9ZAfjiNucyBwPOKGU9Fg9+G0ZeYWXy8//lwdRtmJv6KeHIRYKUNzWYnDyK8
o0SfXwC7kkHrFYFY7Imz2IVQUmH6B4v4K5+g6hPqW9lcCksYaZ8rU5z5xjKOOK+8A8pdtwt2fv+B
9z9fJYqZNsiPiauAj++0skwvIVhuy48FUfBWPxbglvu1IzbOridLFl0K0dSjPc8AUqoFCelbxgt3
nwVe4I0Zhzdp7aV0N+NZ2QPyD6/ZdPD9zxVuYSuRhQ1r1wG91oeZ/7sWZKEdfXLZAwerAFrFAw/h
ZLygpyYFqTA89jw1p5fhwGIL9Pu7ClHpbqt+b7poOINVsJAvjki9zfget8NDFJr+jd5OqGS3iymg
YGA6S5Cw9JaYU159RT8fG+6fDc5at91/l+hENmkEm8MDkRdzvYwlkoN+eVjzi/TYXf+KEJ4GKGsq
nsAExG6RTpMhUAMzbsHY/+1eti5ZKJx0jS80A9MjFrakNL5zXKwhOWzv4DTNQjQXnGuW8uSRkql8
R9qxmhOvvZw9QEC83E52h7oEiCUb8eD05gXzcmNj5avIOzSJmoVtn6msMgbQdkajyhjkb/pXxu2D
vJW2h3a1UAnhvz986FMLrUNNQzKeDiLjqVfUmqjbHyQIZH+BeXI07m0gC5N+XP1OPy/BpgrFsfln
Xn+IL2qVgQXxZo+DiUKxRqt5+nE5FI7cGM+KqwsVnYCo1wlLGI728wYHy/2tKDJ1AxqYVM+LK5Fn
3EKZifNH8IBNkWg8B1V1raFhgfUTAiO99xXq/NB5cknWQupefOqCRJXfErRxTr6wTdGJvhkAVM07
ksfZZrKMGgyfUOKznw5a1lgyWbjHKBuvVyCrlFmiYIdo2uKTqq44Rw0G3eD3uysVwewq33hF72OH
hlMIKzziTlyxPkO7sMSnulzvpXY9FBUnzQ9X8UlMv+L4CPcFIaFmuVKpQ7zGLbwbQZaMBdZFz1CW
Wqy9GBS4b0R64qIq3vcQS87Yb8/HoMDM4TOjz2AeCwESkJXJFQiqNMpOErVp7VQ7DwCF6Ms/NoOt
tzMuuZN+ImHKOpkQaWgM9N/QPGv6KVZ7zFtKs4GMAbw/e+tHJOyHUFyxTJUGhPhTi6AorYH8bWqB
+vDdJb2c4GpcnLIpD/6Y3xthyBwgsUM1jeQlWwIAv2qPY9tanCr8eFfqG6HEjdZygcJE1kSHj0GW
NxKopkaS48p46ABJJRzkahV8Fp8Pqe5voLUPIS1CW1ZqLh3tCmcRVVKHaTCBRTVdAiX+rSWtAkI3
f0YKUUnzFWtiNqk91WllW3KQd0/psng+H2XlR2rRCZ618/IrNW52UYhrdmeJ2XqJZpirsuManVEW
9I2o0jOdBtborHw7CJ1VK/CZlr37dQbZ8hBMn9iTItMZNm/XAQGmRYgx5zk56CULPuT8M6KbIVul
+EUizN938VxAFtH27eCE3vM8OR0IL/oR61M/MzzUrgj+76LqckEZh8NOj/1TW96IS1l+bcFdQJaO
nlGgEztJvNY8EyTkBZWJgGIiDGiJ9H1rmUOMNNzS6g2lj0OIcISHYNSbmQ1EVWIeLYXIxOzUe4gF
nxca9zxdU1HmF8lIpeCaJxapvuW7PHamHTo2oJuG4w7KDuyGuIYWPVcSMFmNX+jd0prVNyTKniGz
3hPRPNrU+aynsd50mycp9T860F1vFmFJyzQcmO6o7iXTod2++WstOF/K28f8vm+oVY/2hUNr6cOj
JgMCDhxdA5fVgqdcgEdLgDPIqAPdHnWNIbIkPn+yXxK7BfNfaVi1x1Xezj/juiVuQX7Wc6x7K/OZ
DTjrh7ArjRmlJFqpsOZtm4WM4YFSUccIz0PNcSTnYgpRIEb5LXZnuAQ78ZINoY3cWamAL/Yk0YFb
7xq0BpAQ+mw907cyHu6p+m5pAIpO6NNJfT/OK6T7RIuKjqJZxSWtAcz9s9COhFjUStsvurQ+CMrY
vC3gkLAgniQP/7axAx92tVyrCj/Xaf4MwBijoRYu2QXPAtF4h+LNxIM682G4HraPHBbdW01loww4
5sT53mzzFrtPTO6JAKlTaPfPV/J1+wNS2KnKFq1fm+hOmiBQaG9ZTQJY2/1U5zqX+5eq2dniroOq
5pIh0wRy3Q2p8c5ElgXioxx362dPva0ebt+tGHC0IhzwhvfucKAQBgb30gjhNm3nqqhHHR13mGFP
LFKZ+5Vgee4XftyF2h9lMI2/KHzY5JweDXiLkUACkwm5epYmLTx8KWZSYxZxbiaI1bHHL+vgUu5T
SVRlrHke07BhwMStUcPgQidSvmqUARG+2+o+9F2oTh0KulvhqPGIAhnJHOmS91Qy72WHol4EZPOD
kV1rGl9swI6vV1fx/p8REWZ9EUmwABowL7+c1Faqe+iIirIFKDLmXRVOiaqQX0/ogFhzSvO3hCb+
V6Q8rhMKHr0dK4s9QMgn8tUgbONFyCeNjlS2UzZgRpYsu6vILW59R9YAJ5lUcpLH2i8QXa/5398l
74cROmO2JbI88jPo4r+0IhmWaA3C5s2Aqid6LFBEDMQ6lhUJmAsA48PZMIIy4Kgm0TUl5KlWHyQp
HyBw1WsGB9SmCmFSev9LwvD9LQMAUo+FLzGOmCRyxesG6zM1SnoinsMLIvkVpmhuz8CTTDx9ffsU
nJEL8lVWHy/pjwIou7piudNT+GUBaoLrwS7/NswRlX66xWvyfxt+2jC1cRXaOe3p9fpxwHQeNvEK
/50O598nPEsp/9txqthCj7oXgBXHylO6S8ikuj2wvJRWdcxRR/IM1vWNdL6aVBu3QaqPSyAecHMi
2+UB5ZwXZGU8P9MXP5hrqD5NEicnDMEUrXfdWSZ/8+p/VNjI+QUu940fEta18th78YrGosdYXv7n
qsTaBK3/+BSjj0MFaW6emr+SCHRweteGiIZe687CSzXrOh2WoiWg8Y0Hi4aRba0PnLNq3IqmnvZ6
i4OqOB1+fyOMeRWX7WZHxD+Z2Eku2wHAFc8ALCgLhizb1nWMdgTQMuiM3LsCJ2OtqQ+F28EjpEQk
EoAOIq0nGOBAVMYpzCe+nSmusYEJFtmRi2pr+yaA63SYVeQdtkObusSdLVBZkgR2nNFQQHhcHcmF
LOVOu7Zu0QXlpKH3La6mGMfUnv3zBgQaPfiL8p/I9r8m5d+aGdDjMbb3VHoqZkcvaZuB7aKcpG1Y
5Fu/zq4RKOV6DAKY27SfqtGgLo77hkVad7mO/5mqi7PRpc57puMEU9qx+OR2MywUY0ExG5nhoTwL
78tK87au7zGAihU7H+RLjYPDRGR22R+up0CXAUE9sMzdhY+4fpGmBA95YB+/6/7PEhmtECpISkij
bOz9TF6mbrkKrspiXiVeGnihaao/43H2RbZR/V1MWeY2hWFizRURDbd63pUXRClCYC9mAConQUOA
hrJlM36aZUiEJLf8nQ81F3rxyk66b/3a378lSOywsqML1QZQOHwkAQXWR+NUv1ukgwlA+nrME5T4
OoAvRbDrS2wXHq2P2z2Biiv3SE5qVpAoXpg9vzUySU3NZSKAXfdrIGkXyhRpVJ+Y24mOZLutq6Ki
Yo/QeaMNXmL3MPVGTLiTl22St+i28JAmDZQdZY4h4/VJh/SuitoxhMkvGb99pc4YjuqW/PEDif4L
7Ml+RAAMuM6lk682YnOqfE/90vdrA8F7Rjwg/HLlk18g+YK0oN8UXw+dVWWjC90+B0umnVySazfe
bCwopRCrY0BvUZ4vyWvnm+x1DzCvCJ7WTAJr9WVAF8tGM5DL0mEgCOcaDPAb64thVZ8QbfL5BO78
D7ELFKUUIYIC/zWCyjP1q2DStCNZMk1YzsqaR+fmrS5cq8htHMLQFp4phZczKWWsLnfSMscGF62O
PtPQqbQ6AT3AVhApPMgVeqHc0TRqnNP1LGdS0OwpzHkbQ5kqSqD4AjTqoavufbGE957IulpATPUy
yITZPcu280Dux/QY3ReG4G4zR3s3tEIWsVeAVnvQ9+8bPKHmrWJ8JuwzJzP7WYDXKoLCciCSOJ/D
rfwJz0i2hsWjG6jUJOBHjimtVgK9EFGVd0UlrShKLWj4XNsU/ukXA9LmEnunTxPJeGXTerRJkKO1
ndTFR6IUjXnSvv4YVSZGzmFuO9Zy0vS24dBYncAe4XzoLwGdPEt/Rg99jgrkbVC5hvA0PC/BvwFc
saQ36A85cjJV4A9x8Y1ukFoPtu1DYmI0PgkLoyQ4IlBl90H+5CjnH2bMWxfHbfGHipY1SkQJCNJU
aa13OPrkpU5eJG4punTehAwywy0j3oXDi6xf8paWbo7T8fh/nSuTIFWou3/Z2glovskOzE/rvyBR
axRLPGfh9GfGtAPEEume5nLigrDSA0IJf2h1o0HqdcUbmmReCyZaH4hhfdbIoLqw7WnFhQUubFKi
p6kzJA2jXnGD653n9eWSLSHwsEwdPcAo06EDl1giEEtpDebYRds44ArB9EBdoNd+8jBUHqimd805
3k+QsUnKuo5hBVI9l1rXMcbz+PcbEsNEWYC5k2qtUerykMOu9GgYxuArSNGzWT3STDIyBgLqOXcc
dmJej8hAAMqcjosMl178pWMJ47e98ptdQWUatR8xxsl2AQ5fcia+KLjq+tTe78NmRqrgXAhWBnSm
jmMyEeDU7MRt1JmSgIPUpUg1nOiS2QdVEIUXJt2P6NVEMz9riyD0FmtmtRVTheQbbPZFd4bOS3+c
sFOfm7Xd3TkNg0ahHfUKG7+GEVrGamuyOckDRWgDYn0Aws/L9QqmOviVv7psjb47c8NXw1oFL8GX
WE8EqUmyleb4Qq6blntzWeNetyUMvCAx7IGUf/p4jx8Kqk2i0YAwm00lRqjyy/1mIxU13OcKH4HP
cpyjB0mehL8iPdgPFOV7gaZ6iJDTrGf6W8NbVaPzIdOfsat/NP0nZpNRnyT5ha+TMSE/Mu5JC8V7
Q+WhR2yOWp4BqCDCkv2AIyAVmeJNwSd2jB4gPXLoO3JYsjeZ1XrxVNVArR5JpItqnDRRhm8VowvF
YWn/zpNiZRTFVEw4gE9eaVLBe3AgAS7ykfNl/8nZSCFgaPjjIqDO8za85YPHSCHJXQCzRDli8rba
qwnIpfgHeVQF4tkFCnKKY+tQG3M4p+SaHDJ1woorig8Lfe8BcHJDFcPF8TK2aII0zrKb6gSlychR
fpw/8E+ESOtvk1bjypDeYwus4+m/B61Zr8wHA4IjoSr8BPzeXqqtVKJIurEw/SMzBAgGfce9XagS
5i93lZqP2iKHp5EnamuVJAO/VG3YHDkOFUf/Nn6ZlA5PvGNImcnDlrMfMwG5E4IItDVpZ6z2QyIu
zHupyTRCuy04vvFY6XlrJNotdhUcStsUa4FZJ66O275IrHeLQhG3yWf2bLJJ/tpiOEH/Yw6+r6a4
5N7RWGO4wO+iPqtIW5MXO//IBDGGdHNgW0+v85pCByunibauFfK+njgy64vjxMyUdRBxWq1nLIOt
DIibTdpg2YeYL1pVvR5Mbg7DhBo9MFKMBl+Z0r9l54cdkhsszLhAF2Srp0TjF/+Ug7eZ+WvriRtf
lLcMyCZWHa0bV9wMEv9RyBtLQ9yrYzcolQbnmTuspKSsPxQDKG2JbAHkX+jrwF1HwC64bciURSHw
WaFQxtc8PV1amDA0sm5ImJq2fF3u51pY8MgAo3itHmefjr89Pn3O0Segvj7RDA8g7ug8Lh55M5Bp
6dx07XkZmJpO5PX04J0RJVbq3wSQB55IPyhH9YdM4GcLztt2fKDHADCYf7xA8I1ZdBjPcIgmYb+3
vRrfndEzoAc5Je+oZsq6jRDpVUf+muQ+k4yAuKCCeR+owLMd/36JbIxH/GrNUMiCq8wM4OvvVis+
pz4wR9NQy8JJal1LJjxOOA51NTa9STL/pI+NIePrh7hTFp7A8aYLHn1uuYaBOG2+hgC25B3chutt
NiFZEuq+M+zlS61naA/wED/uGp0blXJhgKrzQeXM+8iKbeKTIwa68sV3KJ66RGD9wiNv8qGba+Rj
JWxa+UijEqCudOl/mq+xhRUW7+5JoBBSOd92kvuQAGeZPYGYxj6UcgGpknEIK0bV6JylYb72OhH8
68FibWui8C0LD0PFehH0kQ7LL4JVRqkNA4ltnbZHDec8jkyrk7QpEr7ved9Viuid08/kOs+Lo3tJ
MwpskSEddBRQAZJ+HAF0DfiFLBWFz/n+Gzp2r+R73NxK8U4JLXJmGLjQgUJODrYZ+HdqtplwAxLD
sFoPgmfkuD030Z/hHeK8yJvtyhP5v2VEEWjLspKPqPlMVV2zXCYumoi0ROZB1wLOwTiF37AbNAJZ
ftFkqlGy8KK5MXA1/+3w7XSxsozl6Eyt7sahwFAr4bwCrkrWS+RMlJ5mEBWypsIm1xyRpkKwLaRa
ThajdaikmM/I9Y3Y22D+e2S6tks8Hb/pigxv9Mdq5uaFtCJRWxMH55YPg27GX9OhjZUDf00zUkFT
poCqRL7Be51SQ8G8gSDX8QAucXkTSq3vZe3ICQ9Mb8/9fbo0u88AsHXWXWBwt4kQd/rwg+lTN6QE
WmwVZl3MTXunB3km+flN7s8XGGtE7/fb4XXaql+mb34+6Pj5C3xzwBHyO9JJAMRbtuhaAuRzBjy7
B8dKaGyqCcJZlkw2YxBvpy4uUfALq5TmXL7zQsvlsR6akhLgshRmhN3rBOWb1NFBV7g8HfYrxx6o
OKoYoPAkcZF7McLWKxZooligukilb4OCLXFq8zkZ9pamUr1pNqaVbILtR+Tn93lNMzbfmNjJCNh4
XcVz64/2hI6A8DSyrO+8NsV0iqcRuI4KYK4nJdIjFcew9ldSIWXdnxDNe1Ky4mditlE8kSvSdTYb
65NEQiwnW9ueF0Hj1RXyh6GvCGjtRTmdXUZ6J0ZH/dAjjVF7ahR4FIbSmkVYUsb06AAXJpjXi3+r
6q8jdA1koMQowozIEADpoF6U7qszS8oJDMkpPpIRgTdBwf6NNJBw3kgR6524Nhaw/sU0pNO33N6y
Qv8H6kxTO8rrGU3T/8SfQVtNYgdX//kuPSTruKR16+BCF3X1vZEKXmf7fvZpjs82dGwQLqxUeEVI
l7yJwWyWZUdM1di+lSU/rzTQCwKWr7JUphK8h45nVwaxMzatlfxSYlsbBWFYzxLjTeibHqo4KEtc
gxpwb5paJZEFPkRjsEFDdTKr0WyvAJIDEc86FEW91FEtO/64e9Jdkb/Wms+EVRwsxywW2ZlQI/5Y
3V0nUp6XAkWdX+4RowJv/tD9Yaj8MFWO8ezyqtsHxDpOS+g1D59Cg5HHabDX5nsNgEHwDct3g4b5
e8Y8/e8jbVepHdqbFMUZ5Fr98DZty7TIZ+lgWBsF7f42oI9OppUJYbZkeNOYM4+aDsRwWJaFI0UW
mfExUSgJZY8Da7z7q/+QnF0HZ2Am3YAh5yOMUR4l+/FSM5gQopr4VJdKJQhOL0A5A1sFqEZngmUl
sYIg735m2bcsYwDTOQfYf7kPIX97AEIPEX/YbW39D8YHVlx0pXu7HGcp2WpsrhobLab9BuqlKv2/
M4LexJVIun7CbyrJSvFB48pzGIGJbe0MGQbC7bmmyQH3LsIy1RF9szEu+Pz6NbFVsksUl2j+loss
46N8y52ADNi8rvw2ry+hii2BV6qMGqqLo53t5I76/cBfwXsZMvms5MFCwW5IT/9Qp/rZ7ziaRkpO
yAj5tUMkd8VbBN9h/DBI6mOdlr5bg67+YzzmQ14QJCxtgpzR9EAwLgssnbjKLkziONdOaevnW2nl
MqZf4FGqfA9Tpg03DGFNXbXcvmPcIkwCTheYn/Ek96vrZ12EJ/FAhvRYsvAwjDeXpEbURdTqNctt
SDBChUKUFYU+2FysjTWBx5Hm2vJJm45Hmhsxh+P9yYX0gZ3yuuu1oaZGQr34h3yZnUq8ARrSRVgI
7n8qL+p7e1HC5K/vjrrk1RgfpnupPyEypFg9wXZK8Pa7Q9VUaXUQ076coIR2TSiqaF+XxQrCsM+f
LNl34j/iNPa4q4ULKWRCVlNEEQ8dgBz4EsOzq5KfHA3jzWd3KLKEwkX3hZdaEX840isKRz4zP/nA
fNodOJ21KjWR/YX9/PAGmRoWU7Heoj/O3PvPl+AjhEbygRxCHLAbo3Kjovr7oBxbkFE79HO/9l0d
6NoIG2GUUVTUVl358tleYsupsnLHbbi49C152GfG+We7nu3xnoLbtwgtUprorLtZ5RPJG4DRjCVi
rgkiNGt7w51yZDjgcINep24ln6TSETVCf+AYuGwO46uEvYSY3ul7sIoVSvV0JbY0BVFe3bbC0rLw
rCK5SV5oHdFlgkX15SfxFnxHnf1ib4SVI4JoMQd5StK5L1YtCd/fDpA/7eK+GJ62OqFl7Hl2i6Lo
Pf/+dymZgWKWg/6OwsfvsSk+3rT7Ip7maMnp7Jjav35O5rF8taey+iC63/aCJbTvjRu02XXMwTT9
YeEz3fip9o1N+5zChRlskIIxize1Z65v7zQuibvnmpRkDuqnbp96i05HTIumP4SQDSdcgHG7sCbp
p1832FsNC3eywPxWfwwKwq3lz982whkcz8q7Ibz6B4elKGOtM3yAVa1LtH5Jir4a/pdOm8zgJSj9
cRK02hkI2lw1mHOh1VO5OYZYS769W6ByZjU/LKHplSiKX/f8wdCe0i8i73fNhZT3+bviDJLX/o6T
zDGc4YeRheTeNjAOZ2Reya3qSNC9jKkq425vskQ+JI3M8zmEVQKR+/D3R5Hu9a5Thk0dOJ2/8aER
JrBB8/HS34CYvpfLSWdMkoHizSwjyXz1qNRODZfA2tSeOge9cFFcnS0ygBA9ytwBFs4SvksRSIIx
lzktARltQIUS02AJt9bJShQu3KqZTrSVUJOgPDdml+0AkEWx4sXEwqofxA+HbpmPUk7JqAbARjHn
zKt+sLKMpRfXJBhATxbJRhwh+v54yQMTvSfNXfIB04rzYRntv6oKHoAm8xK9K1atNXtfkCd8ylU4
Im0c8leD3b4eVR3ZQqLO1ibhvB3/8d+vEgRxu+smzjSs8+YjKegPw4jeS4/tZuBDndxPn4/dhzuV
8+Qt7C7tYrAW8nxuafaTdVzuKK/XaKot67GGVmCPvJoZbLJCSKxLKbCjAbaTWe3ZI33yk/guFQjd
uHQAv+1NiIsfIfKsancisHwnU7OCH8XvueQ7Da0GLmwEE0XHeOjHmsNB0GIbWrvmX/9cugdhmoxc
dLp5sZE5DdgZW6tbgpBby+aOullmposYAK0We/w+rdEh1VwKtmNYiZ39GMLNC3ykcmcn7NyuImrZ
l8JzjjHWOdItp3Cf3jUPsxPuKieL9pNeIpLcpfUyAWWhgSwl/iTYD+ANw2e/BB1RXRUlndzNMwO2
IEIHwUwNmJYOyRRma14Ez7gHSBNV7cm2c0LKt/BI3jkYAJU2J1iVLit5KwmDP8DzuMzrIe6TKi2D
/TjW9XvQXeDkOXtdB9qMc1ZOETVfY4Pj7nrHJdHvf7NAusKgr6eZF7Gj6lszs8PUmS/0GGSXYdMd
fw8hWU0CLQxl7UoyVKcAUR6vnGWOqZNtkTh9Im+srff1+6BFyRsJkk+AyT6uTAPFlxR2MhRukiRd
V+ce2RIzXBtUkmT4GtRJDgqUV/dYZtyqJUkeQJSqRO14oVxGxdJUzT2yQ6Jx9fQLiKy26y6T65HF
bm/aDY1KZxi3snEZaUCxGyEKfxlUecq5zbMpG0SNP/zUyUVF3WGZ3JBisEkdaxaxs88DunwB2HH5
BW43hSnZB6ZrRQiUbS73SOU53SrUSY6yUHdD7VjRdf0LYF5eswQd/gVcmQQE+ZbSSflaWzQjR9BF
BxZSRGXtKEnT6/FTAUR219dkED5ehswD2BwTdcITQIEp75Jx4er4H1hSbii7CDOSCSVwdG//N3KJ
9ukxM6QrGDbwT4lbVZTJBtUIaK117CK0aJJ4nJwBmKCshnRWfKEppuMmOy0p+zQEK0TbU6v3NiJg
1bYjVmXY2PzIGCxpSYnqB6oCMTrigXltRnZAHBlHbIzxjkebjtaP7oIxup0ZLzdZtkWrHM1GS+ny
44d6OvaB8rQXLDkGIxRpxrkY94cwVWPh/JcYTM/NzMqjn8uwrTKqBOi7HNGXM3UP/x746vfP7qpU
RjcSVxqO0+wBRHDswHRtasAnbIvtH2UZ0vE1m8hkZ57Vz5LowUnZuNpu6UZmGUKYbrG0sQH1cTt1
3naAuIsc4k3xQwHTYaeXd+1N2EYLyJk5q1MhvDm0F2kABERv7wkMXXTVcQpUgxBmdq+0gCP91YPL
IZVzt06dxA4EVQXqTRaFYVrVcZS8OvHbwmCwGWNOjKPU+27Qykqo8M2U/Z4GAjAynwS01YtlgyFW
25qmpuxzve0B6Db0Z1qK6gapmf9XnXaGu/pDaGdlhiw5JzTLhCAyh+rWbfurddZc1BRIigZH+x43
1XvC+FDzG9H65cITBEfLeo9SJdfpDrw9P4kVNpTcKCYboL9x8uNr0fKKCrRexiUfEGKImFAjvXCQ
4PwuF4Yut9EswKZUGtCP1sWia0uJ7dymJK0JcXm8PC42feHp+pZqMORSh9PsNWCuQTUR0pi8+Ry2
3AFiioUHkevMrbReedtl9aIP2iJPY+d6R3mZGnzYogEe9hFtIn4MHkYAsItOh7XlLrCFr60ba1WV
jmGenB5QREVkm1V/1rSuH9feIxWc6kDMN/vvSJlAvxxZ6aqt91Uqs6mxV4NNzx96njPs6KLvN+O2
E/x678/54JngamqXkkk0Uyd2blRhi8Rkkh69H2+wxnqoHDXhZIqObgv7HSK9JSRvl/TAKnIoeZRT
XPN3yPPhwucZHBK1TGiFYqs/c940VQMW4mOVRxJYF8QwRA2btP6vYblOuleHy2tIrkl68hSRSRtQ
K6GKzpckRSOgAjiMd3gQnVzy731xinbLG4xY3++z6iYvUyBG2HImbPPy1zom9Qx7XLWGmFQdVZCE
qhic8qRtv9cnkzFzdyxp9WNSjsFN/GdYsh8zY74tmC3k/eHgYNrM6+YdEyOZSGfHbeVIE8u01QE8
j8Oh0WeE7fbglzXqhDp8DFsT7mXvywusirqrv+1WviEtoXy+OR8fgMMrTwvahadINIAcdLUtwIQu
fLzvPHmyJruXieMkZPEZg/RPwHfRrbjQ7RJWLISMFot9IdMrjxo0WQNTXouVij+/vAnVr43JHXtX
aQGbeIEva+o/B1gxaH0RA5CTzIu6h19IJCYFK0bxFTZzoCLxvIzBdDQkF2IYvk1SmGegv9AhAV/O
PCspecIC9pCSlHBhtf/uIPIhJlZFG0ZjfjoP3oI+enQKuWsGRetH1k8YSAbU7lf8q9Q4vA6jUPUj
QanY5ZVbdQsCHLwOGZgpY7kcl9LzGnw43+0Ag30AgM4saOeyeH1Y8kBJBImqiRFN4oWPVwVC8Xhe
TCTGpeM53c3iLjxX0gxZIamWWb65BnLJpnzUWm60qxwfoJCcEaqaIC8R0+rNh4Mt+1gqOzQ6gJh/
uMqIOD5NrkvuBbjAaEhrEltlJ7jVTh5xJKC3hicLlZ1WjU/nTG3/pz25+yzptL/PWCAliU6cW8T6
Gt8eT9894xI/Uke74fBAWdIcfE0AVuuMWR5OwC7hed28QiN5MZOk4zdkBbtPDek0svT6irygwb4r
rbQ8iZgHJwmY8uqjmDs9nxLLu0MihbxbpbjymspYugq5yHleftf+htl0s2UoW8NtlQv+AtepWhlV
BaeUfeIhQ/2b7QZUT76U/P9I9N9E4G8tuNDiIOh6MRSo7acfDUn8YNcHsA2sxD362CFacZYExSHi
CqTn/X1acbgfhzFVAq69Dyaq3haguGuD9N2ayBO0o1z4M1ptnU7YuUTjFBiJztCXlaQOMWhfCGal
y4PTcGEzuW9j2bTtWfYO8YxQVDImKpf1h9WKMb0RameVuGLUnTgWydvmSucsnHBU9zyVC8sPhqn/
qN7U+F/dpSkPAd2XguM33KIbegxheORJJun3P0mb/go09Tg+Ky2tDw6duw+87zwJ2wDoqlgjpWYZ
Zb1BsUvr+vokDEYFkjjm6QGOWqRjU3L3kQaNlwOr73x7PxkgBtsiQW6TThSuDplsMViGDjpl92af
iBYRZ9fjIFwj/KYrYFQh4qGHolc2qgcVN067BuL6Q1fRVgXcOspWW0PignWsG1X/dNCqxKTZBsoX
FQ9gBOUsvuKfBtq5x9hbcCQLW7OFCtWOOs3h2HPkwyPfXGcdgr7ZY2L9rhJ07JL44N08hOU2hxH6
ckrXm4xJhkvSLWCo3NNX4UD8TGCskwVVEf//TSrxpLxdwiNeSeoIEbpjti1BsB2L1B8mnFkfs0GF
gr5lwhVrqAktWmDe1htRr3/Jiw5YQvmz5G3geBR5zheeIFKxIahSKsF/TVWdBEzktUa6xAIOwbNf
G6J3AvAmB5UkKrSd9wc2tXABkI5ZcGjN8RHTcwS1L+mwKxrJYgUt+u72JZ3BoU4HSnXgrj1bigTf
IhOULc9TzJaXALU8z2H6dJQkSIBUt/+5hTN4ZumKkTUNRDlwvQnmbpkQnIbytlbmsVQWMfo8mjZA
Nb5V9yB0oZzPyhM2sFhd73MYYr77zLhFUHqW/4jOOCdwqtzUb/XsfCSCFwMk7ioJrqhs+ztd3MIX
yH66Q0PG3sxbmKKkIapsiY3PAVokE8k3R4ElV7EwpNZRXsyA+d35Sv1Q7+WYdmw4tjvpYts/tgwo
KmAbyBG82V0Wycu9hOnX790WRZaUfudCTUURvU08n5KvDVloM5DJBQRI9j525MUnJHRCDa+vKusC
uK25+gCdVuemL38jRJOhd18+eFr/RjN8/5J3l1vmCSWIfT+O/5z5Wq2EKTN8kxLWFlRv3g19OIK1
UP4D9VkKbVnZWf9IyfsgRnLc+QJ6Yy/NOEk3RwDaCH0vDoC5D5taDqJHHle4AUKBzuuE1pmHi38l
IvxIR1z8wSBx9o2GDyrT6teGZSI0Sy2ZfF5pwZpaI44mkYqPSHF8UbXdhi0vY3nNiegkRtChACVm
ie4J0hMPodwQjbCgyAN7A1z05oB20RCF1j5C/0hyI2RaHN03uBP8Hxy/LAjm5zwXpYWLGGw9w2Qw
v8WJYHEx4/4+6MJK82lIgs+4Shntwg8E3yIhs0jLMfOnHDPZGcJDQdgmPQm3BSxRJgEU7/2ZUp4e
2CLaZCLKlGYdZp9fMaDRcqGPUMt8wGz9mMHLMtECzwjSh/VyRKgiGo5wUK0/45b0URv63G9zcGOI
DKBA40wKq6y5ClV8oNgmYAZzQNcQP3r1fx9DYEz5rw9Q6aFdR8lDFHlcrMlbFX5UvuCV7zecnfqP
tOqOvThuursdxZ2maeY2scmmvKwlsepxp7V4wacdZGHhYcd30NvsUVotyWO1svrAUcJHnCISIOg8
d3YAtF0embMJ1flUNMetiy5sFcFu/aU5+sNBiTNnvYtYtKGNBTKCENhc9n7iTY/8eJdsyZNlKfEF
Fqb/Re1SXpq9fdq6AAlNqgvuQpQR1YakQnLbDOslVhSd0bxKm732Wyquiko4fOjYuIPd+Yg3THZi
3H0w0b51kp4LjV7BY/bNCqNHenKQVcud3oTNDi7+kBgKRKiIQfV0bVCNRlRpDfSNNJv+hzkxiTBl
89DKZgrsx76ObNI+12F+R448z/NACKnRMEaQkftGDLligPnFwkt6y6dyzXbwSXBfJ5TNQXmbpUPR
2mimge5N9GOhvXMI74kAza+sBZVqa6jkFCs0MT3AiYCezriWB4YVF2UzUgc7EN18QFtJatTZpd4q
lRlxG/rEXOvCM7LA7hABd9P1pJIdfXkWw+VCrNFFczlHy99UmQjyEmzdK5h+wIOrsU6zNbuTZYEs
g6VxsVO1Du6oqdWiDv3CZMoqmzdErCMLSmdbGEOeMx4Nf8oNgukrVAJjrl+mhWC8R04X/M3HhVoK
nv3o0SAyRfn6NnLW1Yvp3nD9G1RmO/D8/5t03kc0AN13Jicir48dcV1fbzeSP1j2vMnnOSFz9qJP
GwDRJwbOoKVFgTX7peh1O6jklPDMdb3ZcOlRvNJMWlx2rz50JCK5bVejKapGXBRvry4xNZdP2bgi
E4dLCeFwpJjO7g6YRpi696o7JBT8OkmB/5ns6vkir74wu7xJ8NWFoM3Bfdw76HjJ+wiGCUpmEtLa
Hss9cg6nsWUPOEkN0A9s8FvJ1vVke3tkvP+jtfIrcCcYb7dTBtdV/MaY8WYoZKo4z3bSeHt10HtI
C4+XNCkGNksHlmkEDxdxFx5ciL9qGzkDaVb6OkD4Pb2uTPR2QJQ6vnpy7OEId/L+UC2jXCgXNq79
kZ5DFHYF3ZKrhBPKV770IsYM5hgvYilxWdApEpURqu53/vDZFUNbtd/Wrz7/NVbQCTBW/Evm6QZD
NNjQUbJO/rK8ChiGqK5wpY41EizphqZzjRZsUBA49+UETWLkQJ4esaAsGkEegWiAYSyqU/OdXpJs
VHfNzcsTlW2f9aEIeaJiyXrcTp8XtEim9+kE06Ct08HApU2tie6k/axdjqxURIHWhIZevdGNwSjJ
QbTWG8hQGDw18GGvhpezqnCttbzUEGA6UljAXHKkttIImCBaYCtOefXFdO+VocaMpqacPJHYYUoz
8F+O8hXwTV+6SsrV0zTzvEIxKRoDHpdZVcVZG0OaP2K2k+ratBCN7VTwse1Hx8wxISz+bhVfShic
KRS/UkZeDP3B8P3P2j9NMBbttVfRGOKcEAuDRAJwyi36GyqgKaw1U4/Ltis2bNT2BxWiGUwu9RmN
LiXQ1njyv4WZ9p9ORuLN/sMWeXTKIYqoN/IlxSH8zq5xmdffVTf6soTc2t1c4qsK/XzudUMvgGik
qopTQ5Ucj47Sn6ecr2RXgYGCeHtmuOMoInLUUfBEBBewSrXuDPYEUGZvy708QfBnlmbfEZ1Rq+Fo
n8ShrqN9dOPOcXUHX57BECcNnZUCaaznY/aEpSJW6I7/BOPWg/ZZ+Ah3M1VHTm7SBKa31/vaIvyA
s0dt4CZimPLJhd6CROhzTYAVUOvoNORiXN7QWAOXM8HW/cIseIZkI/JELSLFG0Jk9ER5umW9gCMd
ptI6OIfL2wwycrO1xo2+iJolXW7QTael1UI+YIT1pB1Kxnq2yt2tgZ5VZ5ih7SO+7ExYssBU23rl
hMhA9O1DtmeK4x53+CaXywGbDIKCT6L76hqYaG+0CXFvqltyIx7VQv8uS6pnG6oqyFJcWEXb5x9I
wjixt3FImaDbpV0zMQVgdTLHAZuNjlMynhC4JkuluZAUy0dEsJspN5yuwz0C5NNjua0tEjOAaGS1
x+08ceU3vP71FEb6bQFgCNBEEPY3Sz7fWPf1rgGl3eDQpzc4IP7M01BJAhcbO3CdE7jIRX8NbNKm
Tw3LW3IqaLNC1CtYC1k1RIBERctuH4NkMsRaxOx0BosKJVqUH/KffexjM9d/Vk5tf5yXMxNcRfYR
CpuxEz5pnrX8L6SLkUZDq6PEKBoVzSY9Tus/oUReV4PJAG0iRZPrWvCbTOibP92zIXp+UEAevgAq
SU1E0DVehjWNtotyi/uyQJ82Y+Zq0lQEhxuL9HUnwHn8UJK/uqFrkcaggADJ6q9Z0lJVs0bpONZ1
XB3L7JVy5hPcB19drS5RxHS9dZepysvBaLTtd0WnwlAv7G2V09N/LmGqRP4lUhLUUvkc9l/wWjwI
qIBPGxqIasINTfH5TfWH400eRZFaBOXCGYLiPeXgrli4SSxUu2E5gWReMHMCyC4VDw8cENM7vsrD
Y2Ec3soReQZy/01d9CjQOezGLhP7SOovL176m9OOhWivuyKucjH/gaEw4mqJwDCz4PRcUcFQROuK
ekyZctPGr4zqZpyp83GrHrmXEe0/RWQjRAVLMKJjf6E9G7PfCm94Psw+P6ij1V0rrfgi1zw4YLTF
sv+ePcX7tDS2WHG0RBhLwqp7M5u38LnFYGFq+6vs+A+iyg96HOZsLzAVd5sFbVzeaXN4gf3/2REg
pf1PTjhqmlRj3UpRw2lI+EYyfGIxJvZbJAu0q57kqiCAq8+jFguj7sL3ZqEXFdg1rcYQRqaftdfz
EzYfdV1TvWszrOPctXY0pjQfI6wgFYgcNSAFKRfeM+H5OeTC/YwfaiPelwA76yBhT+OF+CSEkCgX
QBommWGNlxD7VPbIu+59XcY+koHL+Bbuh5d5CvLE+Hrg55z5sY1O3vQJ+YEKToLJhH6QZsIgD4ju
fZgwAMQqQ35AnKL3/e9wADGI4DAhQhnVawBClkSs07AD3cT1FVJC9SpMpZpmhC0FkiEq1/jdUTOs
nzZe7qkTKWCv5GLqFROMPtuCeg/Hrp8MG0oM4JJG5NDejCp8clAOycY16Y3SbsH561Pf1yTm1d3E
9pb1GHo+cXyu75ba/xnOEdg/Z7CE3Yn+JV7gEJj9xw==
`protect end_protected
