`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
QhSehXUyDurw7ywCoxZaSldQS2za91f9/wgwqih/MLPlu6Je1FOa24AeGYn1f/7NnJAEj3xGkOZT
4ZBBSyWo5g==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ePcQNXYbvz0PkEWzEW14LYoHrV9+Xqi0EP19Y3Ho4xtge1MYNRoNdRWZhY4PuOybTXw4h4QWxuTN
JwfYfNl6dzM7q1JWWH96cfygwFgUZ/pSJLQJ7gus8cQi5INaQ2Z3jLEydep5ee/rGzjz6lKtma+V
w7D4vl5TlNz2UpE77uQ=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
l/9RsfmjItJCDmDrapIifsZAyHbbDmaou/OSfNqFBxp4TMdgrI+ga/eE5eXnvSG3VDo3iQMreC37
/PXdJPI/7RMpuOkSsG9iyuxKn+kWv1LJWKQzi3Yl/0/JWENDV1GOiuKhi2iTkXEisrxlpyp278DY
LC40ixpjEaGpnACQ8wQ=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Led9GJU3esZ32V/vmLYB9/YRd5J1J4LAr/3+W1uQNOYosjyxlv0aMsNDd4K2YnkYb2vkBpLQiZPP
wmE3RzOfIZDThkpi7jHvQjQs1y2BHVmlrrGUC5vYnrY8wukIQldEcmCIbopelmSl8Xed2so6HnuT
B4sL56XHQTqlm1JwfuGDYK1uILoUoMSkU7gJJHKIGe6h/iIePbYanHh5w3aSWtX7JZZf7/2qq6np
hGljC/UsuVkv9wu4Ibk/FdJLZLfqfGyFJjlKoeTfHDKDzq2RYmBPMpdG/AQLz3yZ8lUCkegbPn0N
pyjmqSpAz6iXkDWOaE0ZOAJuA6ywL17jscSrKg==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QINgZBsr2Mwet1cQCg4HjNLdDGkH6rdOk+I1T/lxnhtsAOHp7a5EO9EAYCa77tYZsc/YfnA7eW0A
MJdTtJ3yEcBG2tyRfBONW8WNR3XYJbnHKxmH79XvGgUy43yU+5Lrsp3HK6Jn9tUGasB87qit+WZT
ILJgdTkDRWg5RJbAlFMHBUh4R+qSFnH7bsw4PGG9xvSvx8Hx5AbdKX+Z1/7X1rnLVkFjXl9WhKhm
bjqMA/9ItQ67vc12+L1TdVry/JrTCYr2DOC2MoVp57LbK+xecjxoIt6J5f7caaH5QFt2WeVQKsC3
UHYaC5KLY+yezHeODibzEZq5KPNuTUNqS2Ckvg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Bw6iPTlzMKeyGEG//+fxXTKB4BlemBAuGitIoX566KRcK9Ip5aKxiMUBEiMEILBnvb3Z+UpaQt8T
+fno/Ny6rB0cGXMuBij7CbfVFqvEeJhU9IeVzaDtXRjW6kTr1eUQ6tyUg0COx7yD75AyRxpiPoWK
eAWvPbr+qWtkm8AZ4XQe7zmDyNRYV+RmRaF6Turc7gMGGffiS+XKN/kZAaG4gSLIQGRCAEF1XTsy
YLtdhL3aP5aGtr8+5wcZCmkP/oHDR00sLOKbscknggg3gXeMmZK1ietdvnVVSVc6mBeMoS+xap7p
NhZnQZ7pCYXG3HTWCxSodTE0AwRlmx3ujmwbJg==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 26688)
`protect data_block
bicdNEw6RfHyU8x97Z6x0TV+ubSX08B/jFpT+v8niUtzuT9h3FbWM3QVCU/HB6kVIbFiSnDQMYfs
wG0rDxzVetdn8vn7ferE0CLrzrRa6XntKPW64l3qlBocCWze6h3cgAGjoZvEGQV3xI9c4H/8AYXz
Ya2fvxemKnP5FGuM8fX87n9rzjih9lzm2UzXJcwpOKZHLfPf9YFblUnC1/6Taxux4GZTst24VVtP
po0fBHRD1OsLRORBws4GqaAkFGGuQ+2GwE2/T22ObSj85GXSopnSt6JUyANRQPEIXJv4jUxWKSHg
mBa61Z50o1H1yQjQ+MclZa2IuVvMUfhsELtdLoY4C8RXO2SW/GXQosA2ULHV0CORHh+P/+wOATGp
fyaYoT8LRAQRFVr/+nKJml2hBtIhkmBI8kfPIOcULggucaNUzTYGuNauFNg3yqW9yQArLKMEC221
opkHn7K/IrW7u5hSY+/4748Fn0BHv1zwOHVEOUFVXabr1CiEs4qFXo9r28Fzqz3NMM6fI9qjwtbs
M6YyRFZILKZ/DhYr4FAL6VJsVywrMsnC8yciMdr0HOY7mwpqzA8j9KGjiE+k8wzSvUcO38+M5Zrp
jUxjbR73f3G9ND77EM9aHwmgzi0elb2VlOTcM0l2qGkrwUA2Z//p9ajZ63BSTdld5yFeof4XAggs
e+4gJ7ASSSzOLtjVS9nT+W/8ifoBPMU62eu/gC0htsVdxTcIyLEelY8zzb1CrGKukWwLCTfD8mL9
oVliUMbVWmbZ9jnrZ2xT7+S/6zSsrSYsEgMj5xlY0Bo2iRooB4UWx7G30C/nIgZwI5Yrbdp5C5tl
wYOuJ+BXsQ3UouDwD5vhlksYfKL/Wih18L79OvWRdxORdhkS14a0MseQJwMVWb9JXdw6PG4Q57qY
h4deFMbfuWt3XFlH6APhpGOTJuBEuMqiipqVJVfZpRgESvD3I3Ze+oWybbVH7LhO3G1Vvy3HcztE
8ah1MVaMQvceOBJMmeNDnGzsNLDm8vD0Y0QIR2nuQpF8CwdQjKk8nUN/qEgqnF4/mvhS8i7qzIKC
SXksnhLwojsJN9x4cPURQEmIxjzr0RDOb80r/h6dB/6cGTp4e9MjJyEXamYoSu2QSBdVFXkYwYLN
pjs7oYsZCmH5oIigVvLqhv63UuipDV8XlPG0oJXIO6vJrM/hHRhpTtsd40KT1V0IGCrEr/gILO/p
rQKWk8F/wZ/PPhJIf+edxfI/m/eQBMMk0LpQizO1Ait862PvgpwQjXaeP9Re2GxaSypwYDtHKtHW
3wFdDezPDMhpd7TVLOyfJNLnSvBvzntahXZ4d2R/X4hhjXvGns7j2Qg6Msf+dSPGrLYrSC9vW4wA
PDFyJ1p2HPpoED8BP6Kj0IINEqwCRKcX0Pu+DqZ8yrO8ZZcwiM2p+Fqzs9kqXVN8pLDdumcZ7ok0
PKgyBPAjoWHQ2PXhPpKDsK3Ig8LXXHLyxJNbmJKhkAb8lbPvhV9n7r6jY3cKvPfWlbJaxUOqiux0
7iNS33n2c39hzHHQxXn+FGV6hi+1WCMQaypfgu76rJf9nhszmtKdiz85TYLdR0qq1ZHT0HPjgxWS
+F1BuZG3XVBOzEp++PprLeETicXl8gD16iLTKkpTaMrYvnjMVOjfkig2G1VXZQepJ/UrmLsTB8XW
T/bpdOjYUEJvmlGfJqeZnZOahuKjQeONC5L39CZNxJ2aZkR8k3Y/0H1dKJqGXucC1XfbixB+MQFP
GoN1IE7/itMzpM9mOvDXmtg6Zz5AmxCuXH9uE6rauJY2L9agMKRcfhgIPzEbcV4I8/k/mLLF+tjN
DH6o3lbzdWaE6WqrpGaaBtIx1EA4kBUdEVbwhYsDgJAeAk2c+2maS1PJvD/J8BUKq6iNMjtgEopY
J4NIA8vEp2J6IwVT64RdcivIZCV0xCWoSecoSV9p4aFoZSiufWaxJHJ90kDtFv8tZ+XEXYX87m9w
2U9dge8tTkg52nRz0EQhNgSV56EXdxcE7dfCTa9tJIeuyjL7N6Xr3sgQrfXN9U8RiBJmrGRZ7Ran
jNcSwfx53eGo70GcDQhCjvVGT00gmTcgDHyUe4fiY8eFyL0VCEdEssNA2bHEWYyX9LasQ6cyknHJ
6Aeux9hGC3Y4+Nb2fIGs8wlyN1pQIf6hNYbRorBrqswpAxNBq8sMrIeHVfz4edujcC1/bO/TdsbB
ceD6KZPEY+AAPdJUgy3sR5lW8Nd6IrwqVqAetaG22xrUCNtq6xuKTYs/2tB6VkD7+WDBYMkzR+U0
P6iUDnMkpb/DWdgQUvkP8ZFAvN4Q0xiTgHrBlviw/tFs5eMVzF1w/CZlPHgd4fhCGevcwtaC9FQk
V8o5i8IsjYwhw4kgoq/U6II67txqPliPtSH6+OErAWg0MkEti4zt/d+vmtRuDHrrF1u1RadvvcS6
nKNV+LZ6387E+SwoaC/yGZspO1D+9wXAloysW0g6hFUFmGuQvqVHUq4ATx5ehb5y+Sr9VTY/79D+
wFch/9+qW7PpT1aYQz5jrnzSODezBtEiYqYtniUnbxMO5Pw/NmduPZi7ajGUuwBQpS2gUV14vTi8
zigc5aekK2llQ+INbXlppHwxBLHx8wFMafn6nOgKzcZmfOZCcQ2kY+Yc83aCl2bYG4778YOKFzUo
0c3YOjsy5BZhRPrwAiMzKtQKBatZI1QTQBIND0wfzwEPZOXvtvcrRWLtzsKv+XC3Fd9BBIz3RmMu
RvNP+EQf6tMDWNsC91vor0P55Rgd7wK8GTD+4K3tvUn9kWigDfuZFCPgpXBY040pFKM4TkHH5/2a
5fQrVuiP0gDel8cAomF8uw1+C2BB1WnwFyUhgoGsaeNVanpYCANGe2FSNMc4uZzAFHbSt/zMi/Uc
gi0P4onYUITuglaLimtoxWiHYdmA7/nWrkEQys167Sqo4DPvN9jo4e93Pz/BiAAzGbg8jUJnPZnd
CGrxlRMC3fYZbn2b+qk3ju7i/u22jkdMc2YEB//TYcdBQDaODEo7kesr+nPbdhIjeZscsUBRlDpN
TLe7hH0q9OxZvF8FwzK5hjJoal/1kN8XCTmDNbU+30Z36hgnZJj+YLvKAkaX4i9Ie7Z0QEqpMq/C
bgqNa7ay2lPpAxjFmv1ilE/086VplsQ6WpfhlYENIjL/kGcE4Iu5iqK7eNU2WUiPdABB+W17eEBr
g07Nh8ZrjyZkgqzgjAnVJOA4KUvcSXomUAm6piUAmEFZYNLUEDThL0kB//Q7Rr8RjC9f1Ew8PfUQ
s2qH7txuATlLOHyZ3gR3rUKCl8f3QSok4toZ6613UX1gI3GFU08pPwYIrD/Rs5Enk3FW4/MH+9lD
jjqsHwgE8i1NS2fJxNTlLXNMKmFVoX1q5dhXDCl+k2iHT+sTRutFASLc9tvp4PECgIArZZl/L6EC
xOpcUusWnaKNK5Awr5vEfdD55JJrmGQBLF9iD92LSPMWDQQsFJIS56F36JuBylO66wyaqgn9Wp4q
55/Hs5S3zKFyjLOBlvebbrLIxdErhZKf9xBXfNfxmSYqWwxYmVkx2PTmzEpFI7hZTfqN2MqgzgF8
ReT6Mh8eTJRx6e3hIiOQZvj6gdHw8lSplnqvRlpVi4U362gwJAAn9J9um1+cnXz/n8kAfOYAdvkW
QDCJohx5AxcV+TcmJ0t5xEWyvj6iLMmwB46bln3R2TN89HLR/CyAalEsK0h32VZNgOWRe6orT1BF
/V6dLNk4/QESJbumFa5F/eNOhKvgBILYoACWwJkfoX768dzGVAmqa+dCxmf5s1urb2zp4wK0dp+d
coQHOi0dUIw8i+C7Sr+7SMM2YyDQF7X5aZCLxRXU8kV9FsU8SZcPy8NlAPLgb5FVwZslUNSFObV0
0c2WWGmv0X0Kc82xbKPUIA7/pt7snYEnlRzDD6GWStVXrdUAMKyLS01WXEJaX9VA4jwWL9RXWao9
YsqIqfT1mAG4jRm/v9qfcLhJQQDwxBEIMQNKFhfH1yMtK5R6g4D/HeYbti42T7rmkl1mzx5IS0IB
2E8dwTJffsKbQTSWYCkqmAa50m2nz8r6bAf07sAfzoV4A/BIfuy7/cbFhKAl6+fdI5xttueQ09Lk
39IXmzfKu3u5yF6Kbgv00YwpkUMHuLoBQvslAQdeWuHnXvtOXuNI1JP8dTQUT/8tSHRdT2459jLL
ZeDO5DhOTT59x+PVUq0DI1WQUKNxFnW7f4C+23EFJMZ/HUtEp5ku3iTBMObo8kdgdho1pjjcob+8
cQuwFu45VhZ8B7KPVAxzVLupXrXUuJX3BYjRsfav4wL/S0SfTxfghTSCmOd+gA5c+I6o3GTE2o5E
apeHpOKdVx1rOyrNibZySwmTpZjpWssUPaFQHnXmiv0Dq+XvAdbxtQjcerXFaAeadV+R336XNrO+
zL0vhjhI4sFC7SnnZPP8DqXSiDydEnjunNt6pqav9Sye85S1WbxhtYR8iLBML8oBiq+ddBYlqRui
/xdC45NjOorqeGfY5Lzv1qRYzL9H2ZuXnj8Btjr1gdlRbdtMXugoDK3GLf+G2akLLozcusQojuwY
IHmjkObFKsyH9vgXPyWw44wWPL4iRIL15criocbF9ccFy5Z9kYTDm8JST8VCgCDjiZZYXVF9jqPq
5Eq5z60QKXEqKw/bZY+YYYaK0EC8efHtq6oxca6EFsI55GOnXORWg7siZa8TLdwaFijkx7zXBUNi
mJjc9lF2QEvMEXLReGujIcaKf6yvmE//EtIAahC9GF1hFnSFtOTnXRx0skoeOv/yi/MIZBNMG7ar
7fFBYpwiAAPxKTEc55Bjxn4FWfwE/A9Y10+jmmZFdJG+xpFKUlyRBwsa7DSWcraYkQMjJnH0mMSS
7llJxRxx3EtcobFq6323uLmwpzMawosg8xAVsy9btp61uP9/1h4YsAs6t3R+hBGdFOH2ZAHvGvOm
drsd1p5fL6L4J8K42oauIGywzq15IKgREbbSYsMRX1ULAUQBn+vkZ7fPMI15r5jSuKNBZGjktqMv
0DkXxe4x6y/6OzBHJR+R4nWsKzFty7AmTkp268hhBZBUrjtBXEHzBmqUoNSqfQvzPhlDhiwqcllH
OaB5na17vpCtGY5xW6KQW+OwtfYigjw/LxDCtNwVhB5adhRBIKuKe0SC6LBLFFrGInSWmzTMK/2y
rsW4gcHOxtgpkRF/58316WzB9gmjJrklJXQUDO3U4UaV4pFqEkLF4L3EQNeagNWbNpOw74lZARga
r5k/M41D9WoxM32wjZLrC6eDvWPlYxXqgYIWCpmLAZZe+aXCSjNM0ZtmByZvwZANtw9ETqGlHdOP
+JoOcj3a3F0HeYTD7aJpeBC0sbE8dVjp9GjjmbTs7Os/rWTy9qW0U/39z2vOqb1fR0auzEZvcX/B
I95iohlnqagVf3O6UYwV3iaNyP9yoAxiajhl+SfCGRgRy/QN8iKh0bw3DwQKo7mtjEUTPF3tIq38
yf3P87RK52Z9JDVT8TYnAo3sXsqVm1398ji5OzxuAmKXAzaNGCeWoddur6HPE4uEyDOSSqGzdwAh
4wNbeC7kW8QtQMQSM06hhfqOrB7e6+QxQx0DMLpljfmtlHp/48uxas59CdPjJHShIOrgaQ/h3MRW
UR1sHL3PowR02L9N2+UDFra5QSKlTr3S7i4QSL0SSWluEu6TiZg16f45LUChs+5uwSm9s2JYJCvF
FcknZB4ANte6W1gNbRWrL8BGZXInct7Q0U5WdUgVuBFBBauZcupZUW2SGTxjqj89oKPEY3FBmlSw
7m87xIycfvMnQGC5xWeCLdsVMB5yIAEDSY2+W32wrCZDcRNIffLS8vnrbcNMxCxF+RSYtdqvc1r7
yEVhB6gZ6e3qd66XUx9iUJZH7UyO8d35iXEo+MtbqL42K4/pQ9VoUPsPUoL+/EAYbLveCi/Sgt9r
QjjotjVjwrf+j3ZUAXFOQqf+VjIEm6XMyCTpuffCuePU9tyMnnoBws3p70ivoe1c0plqog+B2LpN
JT3m3Ko7suTRnM4opSuNq0njIUeo1tR3/4vvyghtsct9o9N1bwnT9nMe0DCcChnrRQBAeidE1yUJ
qiBEAR1oz3G8uOGyYAFo4bZ08f4yO/Oqjf0nFEh6D0nK4u0GpO0k2ZdFn0CUo02hBXs7j49F/UgZ
DLs9ZFwtwdiaBnQia6RGSQgFbapTXU2JUVT8DgnZegR8nH+OVUwu+LGfOrArvYlnec7aQ7nqxuzZ
Ar4PDc0weN64dLQEPt7Ljk5ARL0vAQllhUVXXoPR3DntB2JdnJ+dZqQAr8FbSUlgPVjkp8RWr8jP
sAl2AI1/UesHs3YsELL61Qw+bXW5e3yPTHOlk1e0l72RlfvPt/t+Flr5bo0l2pUlWegaex9bWIYk
Qak+hz4Pp5F/0gMhp+w2wEEcCTm5Nfi3hXszeLBT2xYJ46UD5qkwmN8GVfV59Xua+0yBUdypo7NS
Ooh2jtsQHdtgufBxO1asczM4theqiwcky12rSQF/Yughxda0nwl0tdXvZF7ZlRRiYDpOmYn4XrnT
rt4WdowLDmdKU68pQZ4big8yRyurQvG1CKta9cqyccdJ6rLJLE7AZYABrqEn7aGjo6m3I/MMKSTt
XxT5bvptPdqlwZ9EOOFIE7lrHRd7/D6NO2Hk8TEOGoqF/L82V53YFH2b81ECCQMo2UuXH1fUiuXW
sBpvbD7v0CwrIRz5XPSmmQez5D1zVmbrr5gTPMmW2DokRghnvsreR8dt+FcSzO5FZvswPXF4k/8Y
ZqYAPGKZSqBzoDvJXTPKS7ruc0MN/3dC4NDF2qyvzfNg03yy5hQ2IcAMVGrEO1J7lP8O4ul4JJmI
3H0Q+AKzxTiUCou8Djt82atYmRkTKd5ZEw9F2dowUimMXTl8FMhn42ZcNXGdH++lX38D2Spj5EDL
DS5+4QU7usCt8pw7aLgpIJ1fyVuAZTzF6kBqBXx6KSeSpvBCO9kRnRfKe1mUSC6MC9UNHSwbLPjx
A5KRHTe2z0qye3Uuy4kCaHfKJGF17v6xmFUMfCGJ3Ks1eKxY8/JmSxicGefUtddoCvA4P3A+uxjX
Axmpl4G4E8uWgJsQ8xABCcR1THS4+/WtvLWyEG2s98M7X+44FtnTr9NNCtOfAy68MilVaOYIapTm
rvXG55YT5tVi12C/d9hiUOgcwSa6IqE3aSl5N+RC3vzO/bbVFLb1w4Z6Yk2cFbS2IFgMn3zZHbu5
u1jbw/S3cWICRdL32r34U+YltXY97rsguPgnmWOHJFR3M40VXqiFPdEYg3SlVuVoDkO9p1vaN9Ju
2jRr6U6f/yN9yc9znOSSXSPnEYTsIUUIfCw7VwV6hchlDmJR8o5ZpaKIzq92vO0rQHD0/4rvo2tF
MfRpxONsim0d9F2BGYtZ8fmRM3uCt07BQ1FKcLCNftuTDK4EwxuVIrNeDmYqADZ3QVpgXtIyLy1C
MmhWZR6RZDwbETqtQcYkUGRICrRbNT//s3j+0VDTXGpgSfaTm+Stgen5QXezE0oXJmnstsV1/sT3
Nfqh2c7Py0SR/QLZp8I0E5CRBm0obJKd0XylkwL53S+XFjsgzWEowZ5yUSneeCG1fp6LWyjRxdvR
v4Tqqt1e5S6SSUyQ/Q5LgCwEJ7sJgYkF/rwRoSCFC+UxXXV+IHLNzRAL0IzRlMKARp+efR6YkPUk
/e7KjlGcaBJg1nOEyb6dCQFuc0V++75YFv8yZm2fEAPlUIJ+O0zagMg6m8U0/y6bdXVv2w2+w+pY
Y7In+xPJ/gRsOClRRosyNR46f+3F7+qabVe1x20PX522rtO1tD8VGSKrJAlohc9XX2v/VJPLtwSz
vIwVXu7DOOi8NheXUpXZuPVFzi5pceXazv+r05W75f8aSBH6HFdvfbE+Jfx3PUQ9D+OoEo9I21vW
1aORPI8MabCSVFND/SB4d1PjyUK5jjtfOlgRXOd+DpdMwWxQydrqY7al1i6pa5Zh5vhsHklFAGll
10HgHV5hm+ZqH1KItTSGyulhw0whhXvRE1nTNJOF6SEXRZCmeY/4wFVSuUWPF3mjya3fRhZ+qzmW
Iq0EYkRGUSKSGyyZGHQnXFlhVre3/cg4F2cRxjspM7K7sRgkXgyvuJOxbJ5RVYyZ2dxwmrCEo10C
SomW/nEUAJYFMNpR+1AbOZHPvQ34+fQEyVU4MhprDTrUlEwJU1DFnBQSQzRCccAG+6hOl7m5Mkio
747gUFETC1zyU+4SbVZYvZVEkU6h2zTzxchXS4tErso70sOCE1mlNhYt19l5YegDsDm3UZBZ/6sL
hJQ7/0FvTrUeISZawobsBMkSWO6veLPYwoWTGX67MCWExUzt0nPfxDNlklmWZktT36ZMLqhXnLKe
oHvydqX6tnw1HGdwFRH6Jw0T7oP/rNcYm25NZXcoyozrc8mV6+XuLpXM//X4IYcsEmQXKvvAiXuD
STmFfAyyv1XrXjJbPj3dMR8V0zj+BbPPr9LuDW7kVna8eImLyqg6OdSaMyQgd45WSBRpX8VvX83V
ys0NFF7Wj9XtC2LrUQIKkhcwW0hHOCovPF9u8MpEU1v5RB1OX5xouQSICJdw/k27aYdADHl9KqTK
FJ9IZ17igceov3Iv1vrPIJJnmhTTlEbmqYktQURNhjuZ+B7IfezgZ4GlsZS4AwXP7QdoLRlxRh8W
3BaruQWG6B9DpIYAUxATVMgHUcJtnU8+/oNmxQUDzyELNYkFycwZI1aSSMThy96AclCiD1GKY0vT
7HloCjKMG5jlAwxAFCfLblzpjP4nXi3NpKjZmk3120gnDEfIbSGqedd9u3wNh1NC3JU6pSSX1KVd
Osv91Q3gq10a6pv4nuqNJDFipn9bun8I8RthNftmWjRRekhT678MHQSPLBVVxcHpNSddH1tAIvuc
owek7JDcWtOIij3ql/K3j9grO9sggQ8gNg1Du1CeTKMDZpUBNd52Jt3/OEdO3KLZdyXY8H+TYfyv
tvT2d85GOAdaOV9xwQZ9F/2BqjMiwyXXM+HxYIssNmgavOJannj8d3APk9NNfIVZbqr0LTO1UxYd
2IsRafAkrx3xu9eqeON3IFKW8oNGt/nQjYqt9lXrkvcM4w2G9GDeYaSSIenQpXq+V7TxLwHMs9oL
Vc3PqKidkKz64d1uZpbA8IrGpW88pwZZhtrj++9op8TqBaH9w+kEvtXcE4bZ5AiVKbL7K22M1iOx
2vPgGcg5LE3cmTuwIDy9kqH8hT3+CTsgOX07SSZk+IWfHV9ee4q77n/5eUppEBJJfpBuweOoID9G
fqh+GQXyxgf47riCemyF1DPEQj0Xy8KvLfT30RZkrsPWIS5/zNIKcAUCZnsZ3YRiyHaS3RuNReim
FZmSRwZIvnsYwuW2CNuESMogZpwsX0nRrveUqeDc5EXz509akW57eryyieA3DU56vwZVASEg+GKJ
8S+gMhoKP9mfayqF30nl/zi6YZspmaTd0dsp413PHWM+yWagM1q/BteUyxrfEtCxO/QkfLDcN2ZZ
sufpB++MjO5UfCMCEN0/OXyvPdUfDQ613KtWNo/NFphnmC9kRlk6HdL+eFXhyYoZldhZObxyGNdm
FD3LQzxFcZsvAVEJNBKTgtxZb4B4A85FRnVFs7vjTgHubKa0sA3Fp2euDvfDakDDIGkk9pFUrd0F
vuvW1U/C7H5Zv+m4eSDskr91QfMHK21PKuSPCWJt9So5ge39ya4ROz6kqT4zon4zpATiVeNXicQ0
yc8qJZTOU6uXPTvfyNtk9O9naHk0j/YRgxuFNRRlV/x1hDas1pRwhgGgnKS14xqrvSqDJy+TPGCA
WWWh2kFzAm5Jj8J9vp1+axfwJQpuNaTWx7mKm1MvzrISkUeikpgDNtg+q30+H9gEwFtxp3noG+Zm
aSoV2v6yPswk2L/d19J9MtfF9VUzDxxC4wtajoE6mf4se+lb0VTZvs+NplpaIDdLKid84d/U48ed
1JLYeJcF+4ng67zsBVd/mJQmAA8nbFJtm9BsDPl6y1aKO0kNm0EV9zTelgpWcMM4yv4kuAgUgOMg
wXNi2bID8WHfUOUSKXIHnYeFMsCcANgpFQreA3Fd61QJeNIWjUEppBnfmLDv5KwkNeA4b8lRBAeF
6bRcaG0+WwQxpB5eziU3Ys6MsLSmjdjwU2uSoAHi2TUE5EhhHdLB+zyP/krkFht2B++RbO78eO69
il1wS8bYQBuwVUDBvMjj46fzYw0bdEgShviz/LizJeiv7KydRlRss32NV4SnQsMhy/D1eIraKMmN
xlwkMfmiXxuj0sJ2eRuEeRj5E4bLKy45QOjoDk09iaJH/ZpIlKyGs4RBoH2kNayZTDq0FttdLgDT
z1Iz+pbUskNHVmu6bxqcdovF5YlJ+XbW+/YYrOtYXeOWhfPjSsG0T9Ray1LO+sMQQRvxrIhxQk27
NjRsy9z03mFgcPj0RBZYlaMsARPry482iaOnNFlhPERImztz8G0oqPc6141pc/9sKveZzueBkjHR
YfKiBsr9SdZUg0EVmWY1b13LadyHexwd1e3zOF4yjCxCeH0/ooW4coPDTEzJX1V0W0E5cQc5LYCq
4FZOiAz9JKTqizFV1sLDhtHLMjzrQKFsU790WDql5tSLcXk/VsaJi/BCJ6O9vtiVKMivPN3loSZX
8tMNRu8Y3nvRkr6V5O4P1cm0RJdbvA4mhcUTRPZivdq4sYBbnkC1d+AArfKxVoLbdPYseYjWuj09
LSGxS6I74+0ZYPBSWL6J5HX82VDqgdsiwqD1yUe7o58mFZoLKUl3DisO6nTL/MeGkrguvbxf0lL2
8hqCSYiJYKB5da5oseOmp8DwfbVLKU12R3o0+HXW+Nm4JpMU3wCdZjbx0Q5s+69S+XTUC8x0+Alg
eAsopsZP8IF4UneCjYISsi3fnYf4wegAW4PClZCpc9F2Xrqyq8vNEU9230GkB1i/GjHn7sQOtaRO
76zGTaHS3i2OreyUBRIYB2ndqnuuoVt2rnHfNY4ZV3S7I7Xwe0LK7H7hgfVzzYM86OLrZ0XR4D0M
8yhzao96O7vbLTWlpLBJqZk05AltI8hNy7qBlJ9l1Q1gwpjwmEjtH68kNOR0V46lu7tALXagkhrM
LC/SsbUgWR6a1V6JwapGgH+sSdKhoscfIsHR83wDaKNGIJV5Yw4El8NG5umVDXJ+TNJPT+psLTeQ
FcE4yT7YIuWFmchb+DE+nTKhVhawoGQuSSkSQ3Ou2kl4lzDoGf6MIEt0ZgeNei5SclC7eU3vMBii
IpVArWvqyPDoHqATqtOy/kRZbHgNaor3x79a+87WygCwvZmvkXkrA6FxuL7PwxdJ0blErl7D562z
A22vJHJBrKA+tnQLeiHcOao3oh/NPda1Vcu5f4Cy7YHitd02NpUy28PodW5j9iCS+ICCjko2whTQ
f7+olEPK+ne3/CJT88Q7AtQqpUlCX9pUfYwCzE6kQA5qnHpwCapc6g1WSBMYAaSIl6kaVPJcByDq
jFy4DUfR7bR2LFqzxHVZZh0xHadfSqIUcoUHK2DHBaokJWixEk/dwqCsbjXNfyiSpAXQN90cOq78
1SR7qRXRzZ0KdUiZcj/P5PNF9Zddgkd5ZXXlprkeYYhJUk/sN2PfslOUC4j6ofuytpXiSH6h6Y5M
nAj2XHzGAHYLxYO3xMMdpoLU/fIOcp6oCR5uW4iGDcPg0rM4qUq5yvz8VgAzvGl3QwPugVsy2prj
cEMMzII2VjVwNVp43jGePjGIUu1VWEWWwWxGMl2pv4UWP9mDqdaXTnZ+zg7KHp0sEU6hMLr0ZL8j
Gd9akocKzJpPq9XuGFlbiskke4HQYvLOn1g1m1RZeEduUSZToDRgguC/Jhr3l2NchBQJjPHxH+Mh
zj3cFCJQQ+KK5+UewVbLpX8pes4gsqjF8RfxlSVkV1dAdh2LnTKzpuqjMb3YCH6JrFfj3Wsw1ynR
ih0BykJcv4NXLNlLXG9J7g7ErCxlQt47VHYty/VGzEnP13Zaf1S0XXmqLK5Rozt1FW1yu7scGxSM
QYRSEHCfLWN6axkOsj+TnCGiNZiKmvnG364ApiVZqBDSrdpcAOaYB8RFcxPw0zR6mfy4zM+OSdjF
Fcqxt7mgbHaKl6n9dUJECBtR0b+IRrwBBy7GP6L0wM/GrYHUgCik0Ce0jPxDQoSxCtKU5SuWs7ux
ytKIdHC84hNnF/fOiJpJ6ruVU+RYuAzpGpqGAxrIMhOoeAc1JCH7+fJEkxhlXoIFYkgjlvGRkVf1
ZhB6pw2TM5EC5qb2QS12e/hhpwyhNoPFyOb7jsT3QMf6dvSKM2eBSzvelL79dAho7hn7rmhcTJmf
5H5BCAu4Hh/aBRhBsplAPGj2QWeqzBdV9vwPYF63co9DFHOxz4Gdri9a6sRR51Fo/PERyPcfiqVo
97yXTzz4x+6SuEsX8lWrhz66aPctp1sE8UVfNdXAI+eh6YcPOQqA+pKU4CT5mIKE+dNgtqoi8VQM
51rGNyzFOFZ/HX2dlr9ycKKVJgzR3Q0I7Tlef+54IujQaNqA7gUFAjuK1bbpghO6MiTh50tuPyOz
Cqej/J6OMCKR8fbk1z3R3rB6p6lidGa0Zy8kSDFNc8AOHVTFeRi1VEwnMdiXlaSK08nGzBsxOPcN
RSRk58bBhZStXiSR9WvPkSCYM7uH8YTPezAPUheEeXYEp7nkhjMbhv8X26Ril79zlBqudxvAq3rQ
n+HIgKhsIZYGs6zGgRFjFfJlNVlP0ENGDJr9LMPsK0T5gnbqMZOYF/E0jvOnpMbJO7JgPC3nhYQU
FlQqvNtNQCqtBAvMFTeSdRGsOoY8WuihORg8lhIntzO2OKo1tVDE5olIZoKNoV+IOXcXByazYQ6V
pQQAGKOhus70iDQnQCYHXNsJFOJKsn/7y1BH1HMkWL8SQYrmImucBAuL2RfKAqUJql769DiQRqNQ
pkPGHG6us8Hf/bdJYToh4zrShAe/PYc0DGhLH2svNLLSezrakPcYSFBo+RjZxrHLbxz6tQr2t+iw
TDCYgo0nH3HS8aHsxqleFRb05oBZOYtlMDTtLyN/P3E6Lj4lrpk+3P4P2RjAkxxVul0+V3A2P/uM
Uet4uY9nfs5SxoS1k/ceN9CWw9GxHi5TRFBoVTCZvBUh5+HoYwOOCdn3M/DyzFp2Rfsg8DW2h083
TT21mX6/BFX16HGBBzN10nDcW/B7UrJUIJfdtdpSNL9wSPlbhJFfVzDLCuCmZ7GRio3C5xRu4hyi
uS2qW3ObbSWUygte4Ez1MwjKTt4dTKEeaNOCoCDrgRVaa20VoABTdOH/ivdkmhYnSIZ7ymfSBFds
r2MJkDPKlBCcluAKM0kxE0mUZL5Z75bjroqcOgyYKbtATK4tiCOLPBNU7wKZKRtqyDnqQjUWr4GU
z5LJfy6Gx4ppjemtlLE9I0wh8equ6H/RYSmbhWz0kz2tr83U2CnPM19NuZMA/YPEIhVBiw83ZGDM
g/EHSMQXJboY4HBYHv3975NVbiNRYOpMgUtAxbHkEBkMx3RnJMeeM9U71POfc5r+LmUCoDBs/JRM
NKGybHhMyAVqIFvOKHDHFluMk1xtd1VOxvUDndURp1u/5hwAyZTejlz3+caQK6gAK74k5Yv32ekJ
4t33FkBPIj5vgx4HABFhDG9yZaYVpMd7Dwq98DkyKD0GWqrryeMmde72aENDFDKjoxUlDhgcb59f
dcszyDVRFdanACwVQQPLU7fJWpAdvOssQQ5nBzm1LdjURu+DpgkAsKOS8EEye8bDi+RG7JBDkVdW
UqA0hUediYrexRMGrq7Po5GQKxhWMGbWZrE2rPqoEgZ31fEaFY2+SuylcXh9QV/G9whOjIt/6Lwj
/bfZ9s3H61VPgtBXYwCh8L24dg+unvVxeYql1JHXMT34YetGw59NhNZwVxL5dMDYApcXAGIhYJlk
QpFMiIGnpS3NQrJVa6Vm7Ub8T0xMFqqbSNRTmMFm2KA8VyAOob1d4jmNB/Sn9/uIghszUn4APdcr
VU1qp3PN+BJJmXcg/+LFwCBAjf/ddGRFt3PPfAh1WQItoyNTvWMdTKAXbN0pZX7VcPAnTpCz2vIc
oHztwaRYO/WUmTHwPS+suTxI1ocPybfoU+k+WVtGvemxEGzVlPzBFq0d4IavkKI8cH36vZYJz04a
d/+U7gjDbmy3yEno/TmWsfEs+WzYPfSZ47nd2lPq2Ysx8gcmBZ5f7u2mbd6/NaeeQSHrKjpVasYT
T0ECieu7p8x66jG6Tk7Q5BP3syC1NunR9u7Nz52N2mHdz/t1el94iHy66hAyZ4L5Zo323UCeASxp
g9GscBZiIG9WFHl8/P1o6vT4GQIQAVu/T6PqHtA76dhl+E4boTTmF5FWflm/DlYDOdZ7oqcV9XaF
1oqKxNrhgpOBOuyDyChnxr5s1vK0+rUEFWz7fQYC8MSfNNbKWchoMnok7FQbfxDGtn5TEA7d1uIO
/aBmlofZJv04qeB+EQle/bQmS+SHRengRdRBAfuqVtuCEi1p+ASOGC3XaNha75pvFljDZXo7HlfB
V+0Pfg/JmbDclLu7Y22IaN+yR+bLkqkc2bqfdZszwoiizqGHVF9TF14Gh4+/vD6WAczIaqPubNj2
9uh2nRBnnUiVk6GFR3xe0NGotDz7FrsZe5QdqpRuRBvtkxm16kW7Dl9JzbvHZqLn1ArcBQJkvkvH
cd6yGwThOd6lliGwC//bDrvBcd9cbUuZ9MQVLiIjOr2GQoTaZGa49pOyy/lRY4wkvM6RotUVH000
56WD+kFdirP13EG1HGvGJ7HUrfMltZi+MDi7osYuXIhWUJHn3DFfyj3zWk1sXbtTaeWyTtPWoayO
Uu5YyEBep6yUbsBPDbYdWZd33/+DOaUrFrrPQ/pF8pSnn2URDa/wxiGD8L9tGZ3XoKnJHKBUp2lg
oaavsWYnrMQfFTLe5yvabj82bhHBxeA878uOWmTiZc/lpjy2FMMUucO5nQI9QkI0JXqrsfDQzv+D
fmcr6RqzUb9sZyL9wLg0X21xXAQzcRJ+V36SPC4qZ0iSS9+MQU5pMXfxWk96m36fD4hHxfY7UJQG
7Cf/4eQaBcdrfogNU8n2dPtTA1RdbLxJ3shEPi1l6h2vBlkrsvDf8fpC5Dnt9MVZVOr7LwYpSQdV
0oA2xXch4KLMLqeB4wG5ZLEcr36VRocSpa2llEYfdfE0Vb6bia4wRWXATppjBi95/yWQzup0s0kx
AXm0vFDfJGcLUICIVoKOfJdVRgQ8jJfJLdE6ygdSx0tvphcrqq7/bh0tUff/MC7XXk1srH/v5hbx
7XSHWC3ZuPjHtLwSJ4EwmTq+eILuX2D2Bv99U9W1+Ox3KkSkU5OLN9OJze7KPmvu/3K9nMhxINzK
MW9yeE0ykPVwMB0WtgCdDq97IaK7+iM+VdPI6R5RabPpMDpofO1VhB/bjN8YO43v3kerXgyvwkxD
220cf2JdNqPkWG5kGI1r5eO/Drz3ILJpmvnZihvLqc6sR0rIrZeOW+AcsHe2lIvitdWLBpjtvYve
+/I99kLonGfD80HpLcP074IITfv0sMUSSJzH56ooha6gMgoW0tfzo0YtLUnDIb/KHw5ILbpX2v8V
KXgfQf4v0nu+ZxaomSOeaYncDuocUx/wosuruP4msfExt25NciEWVzwID0wIDLNsy3Q+WTYYVp+R
/5LpqY2jQJ7MAO/WUWh9BWhfvL6hqGWWFMk1DZUbxaUUed+rrQp9lGkAuNIz1YJmcRKAcDC+dVrA
/Yg2+uUdNd4ttaO4xpMISzLccM7i656hhKiXM6Z3L2OVR/BP1hE7XY91rdtIg0itikC7F4CHTNxD
/LSTM5B2sXuIvNFjIk1x/FDXFoc46QeXDV4gXYN3gGt3R0OdWFvVYTU43ff0Zje3nfufWdAPHD9B
INzG2fntcDinHsi8xNqA6CUNppVddV6S/HQLYzjTxxQdaK7FO0OXWmU67ViRXbM0MtQESeYrZukK
fOVMaIMJHqZfvupLMRI9am8ZM7EEAejJ+cMolr/aLRwFo2UQRx5RxIe5AICCPLtg9tFBNjVEBB/5
yoB5OEnUiDZRhYew3dxuemHYZ3VCejo9OFA0mwmP4HE8dtOeK7525aVLJsqX0reL2UjOgbR96wl1
dU9/m1rCmZx9T36Hw7ynRHeVbxdjuob2h7ahJz0lz+xwJciE5o+qtKy4tu2owIdxO0cAdAv78rmF
fPzNdACg/Kps5OoQ5MBZjGaTvc1TH7qMu1utnMLURGTSZaTmgHPajqmh9VQyILpU2Yog7/OOnNSm
T1d5xItMhuOdfD9B05mng0o3Xydc+KYacdqGUCgOBS9sf3PvjvGtWjzllj3BpsuyAMii+b2BwFls
eJPrGJ/60z8jqpTi5RURuwrwSkIAUXEgdHpbYbIK2+M/z0C2FeQDiO7Hawsn2oT+OAza1VKdnENj
Nx1JUMvRddnIkqN2PX1QNdAZKgYhQT4LAONmCkgK2gS0hu+Qa3FvkG/vsBrqGJJFBfn2dISQNXVc
Xqv7s7Iz/OcghDGokkvKF8CgRisrBveA37ZwcA4np9YeIQOZFZi2jNsHByD/pRI5q4hj/692RVSE
JlB+I1Jq2W3+9IzE+917p6z4YFg59sx743IWFQwDbkXud+2VzCMIeRScuUqXec9tkyGKCiM6o0ZU
xh1AVplmFhK3n0iiPNWGZiqejz9fg3ObTbWp8cdR7zncOVW22Fo95z3viwM3lm2gC+p+o2LQscsl
OKU4KmHEjY4wPkcMtrlEji9RRmPgAqh5ijxfbz9ctXOrDvwqDDEtSoSPW/gKE+aibjlT6BCl4mrv
u9IRRd1g2pPtPyc0n19NcxNnKrHUNd48S2747VOousQ1iWaY5CDEGRldGUyFHG1/dWGqNDa6oiqr
3mmVhF3QM+D+p+c1upZiVjeYsKgx+vfBQvF3j7Rndutvr2oDBT6bgiXZHBZWeb1OeM+Jg1l/FPSm
7b+hOnBP6yQyH8WxepawQNStUXpdJRLOrECCziyUYqxmQ5KVgwd1vNrjRbBdLYMrMYWMgY3TCeHE
tr4qO1ddiK8ePbK6QT0oPK2nDrcD8Gl5Oswdi5KVWBiO/1PzkkZc30zOw9o0XyhdAUJVCPhoorXx
WknpbTjRUQCewVfjHFg+qUIj8Gaulv3VMI3OtLGnrWEmupDZUZzWFi41OFx9l8fBvVVcMQHGprKp
FuA5nXa6sWZGJ2fEozFyU6PGQllIcYeMFJoszJJ94+8PCO2WgfKLT41EJBFFp0JGzHzhBW6r4CSu
8RcE0JEW87DjtaUfSv3AEDdTrlfsPpSU7beOe0/16qZ4f9C+hTwFAr17xz0dNFFOnFBOOJm1tKwC
hN1zu5Rsff9n7wXt0lHVzxvLWyB/5h4D2EvqdyJ/qtPgmTZnzV2sDXklEBTZF3qPnG8OKJqJjNyy
11ZeptZrgEaFD3Plza00Gvj6JfrO3p7k6S+TjaEshV4qIuwJBjMVUGRhjWzdpeyt145JP73KmveA
coFiS4PU3dioN7iU6CTwt0U5vqa6QYgDyd+3QG8yTitr+7iq3ur5XDyhFDaj1K0+SOT2iM0ItlFs
0K4/2D6RG7JnIvx0A/rPIxaITrIW9Azh0KtC1BpuDzrNQcbZ/x33mpNuVLr3AkP3CL+wwYDWpTG5
yhhyceFbInj3MVqwM2Oq8GKcsjYRJn5JzljQifZDD0jbehahVSQnp+q7gvd6GRhb9jwaY7bXZFQC
LoX5kxBvZVx2GZ0DBvh4tIpP/PaJi3StgXzkt/F21OfLtxeQ/OxGKXWLS3HqE3wZvYOuWICEovAY
2jL9nK2AxW9Mah8lzvzrmHn0h85qGSM6VEm9+bfFblMwjAGb55XjUqTn/xRGzDHFefXLHW4zN2ae
88YRl8C22Ei8GobLW19KgJXchnBFa3JaojaxBfgPwb/+MZn7Bi3dxBf3aGeIo5znqoLaVzilMrcn
K4w/q+NRkG1SRyGLNpQM6K/lZlLQJUoVGRP1YDVhp1fbAef2dxFQ+I/gov7ZY6a6eDoF0My/LADs
7f9OUwXSRWzQFbZ56VyBEDAvfTxJYwVJj0mOT0073Pnz15zrUnxx0xIMsgJYN/pEdJIQmtKBoK9V
SLhEd1XzlICQY7EuFVvYgApdhCX6ML+ShRa+thQXeuLAcy0RNLksEYza5qtvohtOoNRNflvdY75m
BX2Nnh7HMKlc+wVBjFffugXS57y5wira0puE7NOKy0IV0wNENFLSU09op6j2hkRO7XQmu2Wh+nhb
3gwyDRGc3pYuczsKTBooKDcJFApRu7gmRNa7oNcXjGxLO8LZZUHYLQHFWetCAViuWqMeVb+GhYpq
6HcnF6DYtakT9lT6qBRsC4bG66dswOyCR733LVza7wr9Mf59ThcMi1cGyoy/ERZrGf5kQReU5Nol
wO/btwkA18jHthPNKzEjwdMfgeEuqXGxHPNSbv6X7b9Gdd3+E3Ux/vcxbGnpq53bx77flXXb0pqD
7t+xeBRc090/IC861cFZisntEQr3mEDC5mL/LqoqCj8bo/G0CLUnU1+i5cEoYRTiHZQLF0LVWayw
TEYvVKBCn/4+4s1795ksMndBV5BfUJIvMKpEIX6sapNG0CP5gL9/RRnxR/pIFarBL78qM5sOoCL5
bO5enhhA+mnaHotKujN4ob6VTwx4lZHlGTl1EwH5EnqhG/2CZplb9469Aod2C0Pgih3Jt6V8nMIW
fzCBHbLvvMnlNGRiVUSOxZ2AZt4IffrIpr/QJLWMJrRlc6bUVyC3KGqUHTsnEM12OdNnwlRnlQxw
oQkkEJcTai4or2J+lhORD80V1UuoKEBpdNFMknsrDvJINZ4vh5DkFZL5oZkF698nj5pJeQIgf579
SS0tKBoyuxqoZdqxQBUEZB/UuBcOG9yxzbPQVnZDhQvi8gjUBI8nF81ix0J1ayIjhZ7dRpOBS1IX
re9Mw4k8t8+T5FEiRzeLsvrlPk0Yw22R/N5V7bydCb6UJ7ClJLlnXJrf0IriU/rUfEuWNjW5GBaK
oVBWYDStVW+jFDHYB17Uy2XdZOCNYJGZoNObJiWO3FgJ1jHZvKp11sHKYKdOqlQlCVavtaWTRyGG
dmvvesqfP8TIF3epNfZrNB2u6+f6iC8p/BVeg6JMHPzKXzZDVNzZBbcMdmmLj+ZtK8xDr0SQQCCS
ugLR3cqWyua7XuRlNT7bocTaw3bfHRKtxnqwRfIw0Ql5nmv5z/U+O9ryZFu76t4sF/IpCjGsE6Wu
nYAzDMShfnONmboKB7MTiHjkEfYtPWHn0Nh+LL1P4cWQwCARYTKhgwbbnu+sWX3ezf/He7MW9Eas
ME/0c8Av1f19a3MK7BLJy15dt3RWSwwTlWJ8bPxuxXKZ9er0Aoz1gTGiTODj4AFvYEANsQ+VqyyC
xdRCJst/oSljsfCm3lskIgJc7w5jMSzOfAukndfSCK/MOTEv/j8X77DC8Y9z/WUQ6ewRBPyxZgez
buIBz2j86XU12cprqrJulUGQlIpfF6i4za3j14tJmv0Njo8fhBC+z0X8rYkJpcgqGwgubLhJPQzT
ZAj0gFX4HXDDltNUh8TwijIOT/FTcH+a9ggDQrWRyWiL4VCmBM8AHtvdHRedY7i7trVazdB7L5gT
iGPiJSp9q6IfxzxH2J0U4HtHV23YPuuDEn9Zbj2KXqyGemRlr2SZpTX2QNUAf8XbmN0CyoZzwzHI
bsXG3dbf9wVp+YLG+AllLRqsLlSle6MzMpU2zV9B6FOy7FpjUN2fYLijugxuUF/ZszMT4tNGzUq/
ijMleODYLCA6d0+aMvnO7rls4A6jyFdNxLoRSZCJtuIkZuPNnf220iqESYPuSfT7yjbE8ZJJmmx4
dKdoHNhzcYh/IzdNtJ6kSYHBb/VC9A6Vwa/1fkipw36ZTHPzbbPCmBir38MuHWCpJ7XuNlgVX1s+
vbyYPmp5hWvN9JxCGpV+Ss0rPub5eu3KQqxvg/7I5ACURsNqBWe8VV+J6Yl+7vIVA35w9xO+z/Te
mWzG69Keaq1McyaEH+Jn//k+pxOYXe3Tu1isn7/w9Gq4XqSKFpAG7rlseYKOB4uv89au25so8RQo
XGnSqQlWdUevlhzzlOgwmO+mguunfV1FyF5PuesFy6WjNQ7OVWFeR4YlWPNI+K61zAKxVwVbZMrn
5m2Wwrf6BPi1aKhElC0Yu14LGQnIppygKZUy7czRXkH1S5oYBlER/6z/somQ4jodl7hMLEQ/bufY
rL5yWm/j4h1Lo6ul8sb3XfGqC54SjUQCjF1kjrExHXRB6ra22lOYwVaDQQfTEFCSgBjAmKIIX0a9
q4eUY/Wf8GxnQQVK5geXw0xP5m+ejUO3TzbAWwraHwfduxfElaqNtltnCMf9d1dZd1bCFXPI21Tk
6e4htipg7tammvbHXtTqo2umehrltPS9rhfJ60Zx5v9GWRQvKWK2452qYFi3clCsKLs3+kOEU3qx
1JRVXZEnjTxeXZUocuo/+od8SCOeKnm2bRkBtSIifWs2VczGeTsjHcdM3lxCUcBcIsqaz8vo8kPZ
/D46HbVRLKuyY57mSqMwihOrxHi8ZNm2cSBV5JgktD8/smfrnxThfNUEpc3gdMmh142gCSXy14EA
reFBRfBmzAEz8d7OQsCNlddsoh8v+xiD5prh6L4DvrqHi5klSe8FUSdZXHK0D2FLEa/liB87CBmD
EZF4GN/QXW1Zdna0jePut6T4hLnHgO5cW7FlD1ABRBIs+i8G8OIjDGjhWQKtPE3TF0jbia2cUg2U
3rvTNE+YbkPMM2PGEi9baYxHsrdEnTLbLii/oFAbGcyzHrPL5XIU4tbKf63T+ysK/iOFs0uA7X+q
jAPgPIa9YcoDrJvL5DdTAeBCT6VGdeRGTSV3quClpr3iB/6Mti1vsrT0oxUVVVdGdIbe/pvecBi0
6do3+gT3Cdrvk2yD4D51x37tpWCM3gvA/P2ULLFWcwBfNxVcVaaQvM8V4FnpTVhM+tL0U6SClJGA
TeqZjIjOZy9L0RhcnAOuw/je6jsrxG+xp1tMU0S2Gw+uV2VrZqUSnvBjsthUWuOHG1sHk+XQ2d+l
utNBYewMNIEk/K5MG7rRlifRPcHWsVMN9FoQCcUjs8SDTqk1LKZst2CT78Fx7Q69+qS5ua05wLhj
Vsx8YeWhSgkyzSEszaAsBrygSxG545IZQgSe8OHDyGVZmlRJ8ECT1oys7RtsO7SaVgTvP/JlIkk0
we9yEGFajdEt18sGgLIElUiOHslzUUX8oCazEoKPZBrWgsSWnsygkqEhiwtCmU/25Tq+5DKYqO4g
1D8NXGo9b/4194oX9Z8laLgGkI4+toUd+0g50daEoGHGr5RIYYq6Sfq2FQ34KBF6G2Je0KWNLZOB
qoOeuddiAIruzgrIEeRype1msTFoNDFuPSPXjEuYXDVotZlxJbVu92eDcuJdMRSgkamc+Ll9Mq0q
j301/iz/Y+sl/v5a21Zmfh99GA3VNRmEeVxS6saYGrrenEEu6WHt9iARNMMP4VtDN3WZGcsKTwV6
iW1rb9HMp52GdfivtimyJmZzbjuX4xjVmF1dJY2wWDimPUZZ8h8H2r2WtFA97pwY1ROouuoeNz57
4K10AAo/Hp+iDTI5dvWRrHoqiSg+bI11aqMcWsPzZGW3HFUDFAcWP5h97xBsWSnFWKFV+31VMtu/
zOSLvWShEvULXSp4BIA4X2CsTkSQjuQi4bISGOuEJStU0TcQcJxMdFpjY6kNsfKO7Y5FJ/b/IRM2
CmhICNfdnMg7vHtq7s6H/Lm4DvFnpHSEnH49cIgI28gBPQi8YfpyM1bodA5hXTohBhezgcl+Y6MY
NRkYjQC74IZe6ADXh37Lyltip40ACC7kd9mkmPIB4QImymxCaicrMESmJPR2OPliKpgLbtmTisZs
vkC839NC6w7l9aVAdTwzRzg1yA5YGVGLc7ThhFM318RGa9Vp4YHDFBdNHmLHvS7hz1BXR0zsYF64
VjrzEkeMQSmGEJKg20knEA7ZccImPegcfNIOtdsCyPCB5/9QIZzbHmowxj+rQ4dMqrb08OGZvJ1a
ziL/1+vcF1gSZ4Kts7iNlneRHzjpPbszZI5r6sg7ZLiOdYbZm7X7otiR9OVlpBtzYxhubmehOd1n
4b36BlTnPxrQhEM6UKe4TkJXYNts6l6qlKDN/tZ1WyoZNocAQngHBCZskM6R/MM5KPaEEQ/ihjJ+
k14Hq2XB92+modW/UQRHU4Ev1ty6bNu0B/4WJ2wA2L4l+W2jt9u67oQe5vGt+/4ehLn9GClSvFjf
PXfDz+70fNE50A7/u7tNBelREfo7Z5locgaKX4l2HaNmpIBoB9zUcTd1MV8vdUIWyNrzi8ToAxqp
e5m8lFUzHxAcsmTYDqoL6n56mqXeBTo443acfaXSUMTg22shrBumyYknhQfdZxNIKPn1w+05O/Cv
G79KiZIWCaUwt7uNUw2mv4ICff+M2qvRP3BklS5pirNQjbhPADaoZn2FGLLYgldVqDcSg8ahBMeA
tuo0cYC5nwmlBCv+db8/fzHyFGN18KBzS5ocEzQ7rw0Bsa9Nq9qY7lEUSJfYgVJJSqe5mVu936xS
w+daA9cj8iR3g4l47KZDh/Ta79xCNraNFj6O+t1sJISA7gy01cEX7fKRczUHrcpwXv6fMkG9rDFq
n6rnPlHOiOKweDIqV1jmYXeZdQlJaNqtUGrcfGvRVY0Wmisxq7qiqsDejmd5L7KcTa2QdmZua0ni
1591adAapKK8Q2X3/tyWSRHJLqJ89HlVOixiOxHRrCUeD80oGZlG79xiXUtT1k8UQHJ9o6BK65Ua
fWElOxmqJQf1TwDwUuGms9XLimAGEc/7dJQjpOirYMW5euUOG12h3C/xl1uzq3o0KlIZ8Cu/RpSF
MFFn7d4GkY1eKjqbd4GHi2MgcnyK9oaPnQCtKQ+yPdL9dGkHirXuPfzSoJPZDPMPC9JNVEhWGVPB
0608DfAhm/69wfQyJSbBYh5LpdxnWI1xaJYaxPai5U9SHC07tfMp2qJDJu/LZKc1u+t5vMsz1rdA
hYaSxGjnN3XLhkwrD0dcIxy2gKkOZO1TyKE3/7i33N6rslFIWh2DpGps8mXnXDxe70X7+J2kKDA+
OvpqhXJJgvr7lvwpDqveO1HRKj3PvU6PZ3J2vgaY3z1n0Bc5jXDhv1D2y1z+BLoQM2l/iWrL3f9X
LhVeL6MnKKWbPSkq4UhT1ex2m8Ymy/lYd8cAbTeEE7V17dwzIpR1PW+IXW5IYN9saSDXpvQ6eVQ1
VGc+Xn9yP2ExurcmxLQQ9rLI2BTFdVIKM/R5olG/qxU8CSZO7uqq6y+q0PvrOnBlwdh2OTs0LaZA
MkjhLD9+W5tHXUQcOzjXE78vsgBMGJRGk84nqP8HqPER+FSvREHOwwue6gx8ndsdtNJUGNekXjLI
aelos4Icr9byUUYLtbHlcxJWZCuukvY1MuToilmKCbuo1g+ky3GBm3Oe8UySolAbfQ7vL5TOjpIQ
IRZgfRM7Q2csHQV8ikW+2bxk2wUAu6sY7PRcku4hpqUxICyEO8swC0RESgTANBuNyrOwnxLsJ31l
Y+7CHTseX1GbuUCTEx8hMvfF/wisLDSBuzkTqPCOnoSBSIuQbJfUr883LfGQOjwwehOOPs0JGikz
lHPiPItHpN+0hQ6J4xzMuxiBdXF/k1yZ6n1c4piSmKSSpFJf0ms7dR4H6k87HtTJyJeh1pP9cwzX
Oj3BG2/gK3qPSR4UUwjrfPdjZxwkDPAHurnad3QNW7g8r+hD5dOZaq7wYTPRXRA1qXxPiaSKlxy7
pGiz/XaHpi368+HFqypruRh6yVWbL2+oKdt1kd8uD8dwD3PH4kKTdX2j7QcsvMm1j5A0gLRLJ5JL
GaY01u2+RyGaTqu3h/Y27dTL0TGmgEVVTCAOBA+CBX+uFYYAUxaatYzB1zhHd3F1+lrMIWK0X75J
IsiFnKhltLBHW4M0BBjzk+oZUYRY2xLV37jdOavNRM0ZxogCjix9fd7Xi9WxmNrJ4aWuvavoFYVf
wVSOPMkqrMkh/g8J5ifZ2s034uJ1A7dlzztzfDQ1LOzaU1Es6fZ0Fx4yT6nLh85CdiutPONKIQPf
kpN2yQuyGYc+Tf6FIRYfRDsqYWkzJyhLUMkM7p0ondBXfZzg2Q0lh18XVEM+MfnRaeCkYdQzj5m9
xEwSHIn3Daqj7IIacY3WXZLckm5WafyFxNtqVNoFPEWB38wQKbsWfEUvB13BPJ2peAu57cAsnggW
qp0rTEuuONwZrphzNVNAlL/8PVkemZgWP7BC1jXvg9uZOx77c7jHQQ3skMt0XT0Hfo0uLvCMGA0X
RajVvQUYmEN/jUgzOqhg6NPm3iMHqax0fUUkZT0Hv48nTQNR6TynXI4jo0M8uMxnzmHHU5IKtTJ4
wha2PVzW/42cYdnLVC2inSvt+mh7bd7GpQRBLI7Yz9/njsxPWkMwyJPa7FtaTkfZ3WD7NeoqaKDb
59+ss3n9qllWjItCIacyAaCUEf792Rpv500VC8o8ih13URzOAWHkUOXs+j6PM8wxvXCzSYtqQCok
wX+48UKsEc/k6/RipmivLQ7xw/Mtd8zqBEdjYdB4cnG6XpswVIRCAVd5UD/KPjLeshv2H2fc2esD
3xNOl7xtQLP6bwa9mlzhxadCZ/tRlintQjPUrY0iwzESTOaTjbx1ih4YZdbklDML6wu4RJk00FfA
bgptzJ2VJ2u2heQS+NktG51I/cCD9sde9ggczJJIShN9VfM1lR0fITvwc40/VqQ4BIJDbLZ9MrUp
tc/ZUgPpaCSYMlYiGFC5TG576pd+5+j4rOhBtpG8QqPWP5ZhT86WhiwgE+p8ztzt6x73G1RKxizX
3g3+oRRiirHyxXF5howaLObhYz8i4Pk/gvhAPygFWFfPqHuJ9K5RqCzmvGqT+IFhnLw+y5fR61U0
94IvzKvRVUU3C4dnRGfeCSfVfsgiXc4dKruD5nzcA7z70LuQDZRM5JsFbpzp2YxWpz4ah4USKu3O
PWgR94uIXd3LBZKho6SJrzvn0Yn2VyIHOSj8rFaps6rLjUEYDu9WJVz4H3zcehUZfrR7Uwyts4aI
EQS6JdpbhN/kWLQREOVMu7ojrBfYkkypnPn8iksbSM5HBEuPz+bTVF1AFH0l10hQegKCof6poRnC
eLYcKb699s5f/6MJeGtCglnhvC22DWXJr/fp0AaWfKwtvP9QlY4TZH25rd8p0P547zseob7lDtJa
2TDErddrRM9/xajE9xoElG3jqJhw8wzPkyOCIujKwTKEN7pyXNsxh6AQ+g2OMQ4DJ5GUF96tMwbV
m/wVTzi/Sw0PknLdTLDqo5CMClhXqw3foolYQ2dcSwfl1ZQ2o4uDlvgzXXw5saKDAWSPNmuk/Dj1
+T33cMrai2Qx3ROLZGhyfl7BIfsOqpOHVp4FfI091gReowRwZT1kHEiOZ3te3CwcjtY05I3FpKtW
7YFVoYFcPiX4kLIYxu5UXF8OnoRnjOXcvzAD73TinWGIHrjf016E0hwrI9F+Kr8v2C3YTlpLabIn
qD1hPxRvKnZPdHIgcRFj6fNQc1ty1wdrzKPYAlPRyZX3iY3IXESRopSn48sWtfeGoK75fT5W+MQj
omswGvFRWkEpYhD3E7boaSWj1P/tUZF0ZFq8oUE5lNJzMXFn2Gls44QOv5hKVMMD8Gkt6LASNSQ9
p4qhzKuiqvCNpZyMxGhxif5PCDncn/QSFD5plcvqMFZwLvvRa9rMQZJDmzPCZYlQ6ezf8H0xObiO
EumvRxjQ0Z6z53BWP39D+wSo+6/LRzXAquUopwWfn70cI2zI2BmWXSJi9GVMJLSTsmWKpi0XHmFa
Rs07IzgpggaMNoPTp7ivXpH/5RGQlAExbmsVAhJ780dXC0ioV6BKD5kV7jnXlnz09TesCn/1VJLY
Bb/iGmusQj3VABW82samM0QcqLjDi0TMBMHVkcR5MMaFByUxDkAth4E+igSy7VsbU5i3LMrum/HF
ZgUXQ2peSAXt6N/t1zNBTDzrUiCkofFpOH+H6w8F67LcMYViqZjBGrFBtfVKj44bwv2E1gTb8s5z
jRj3t0i3bkHB+8xq4fHD+9zxt9JXnbIuIRwV8Pq+ElGG+rq6w32+hNkAzioE13vkjhZsHc7WAaRx
sxgQDkaF6QHw+CKzqvfEGo4EDCoO8+YGOg3XcHgSZDhwDMH5O0qtHyO4kKrfZbQYE+Yt5aogvDhi
o5nl6zpkz5aRUNJr611yIi4C6mznAMXg5vRq+O9zZjhw8gdQeZ0DKLYiZMIT8kcYZFUpf6qbYFkV
Ofz+q636at09EXR89/pz0V3rroNTPUYJ7pVZBiQpd8H3nCz6XHHhkAA4NhsY8JUojnANRbWAle3y
cqfoyWMZmFr86/x15BkOSNakl+IkhKikCWdPHQP928kL7t8lQNMN6zNkdLQFdsdZwpRJTB5+VCFP
bK5st0wx4YxVbp8go9FH9KpHZYB9HeVdxtJQStF4+L3Snay9ZjJ85p8s4b2pfjWhW5f4LVKyylL3
IbO7zhW0yu5MLcU4BKisglkXhkQnKVAilMYcjmkcaIeG3BcQTHBhB3KDqlxBb/dcG1mxEYRODh2X
inBN14N2EWst5cqUJfpM0aQ0xhRf1U2ZrKY+VYZafAvw+Lq9uMZ3PMIheSZ5r0BEJzu1Cr6lE4WK
EErCC7h9PI7yX2N4dsAWYiEdq+qtaJQRBI1sYCBsq8R7Llni2sxc12KzYMCfhVmUy5shjx7pbJej
Wp9GvFoK7RZzldZxSMhDz4+zlfTnYVNHUJfleIczzsdyV6B4YEcvfCQ90kk1vM5WGTURQgxWTuFx
TdLCNQ4qotxcdWu/LxXhxx7DoVVVy2snGUNbNKkN1vvT2tGqCitYE5KCScZ6hKOxpyyoxilVmGLy
J6sfu8DNqwX5B2qTBZfXOT9QXQqB9zEH1BcaBcaIIBNO41Pc7UIrSB2guilCISauZx0cOHh631XQ
8DcWF12QYA0DJKDefYj7Xzism9GkAbNoyk6uGT6LTsXo6CGnTxzHDy7xefY3j2Hih7RarL7ODX/0
9l4VL3Ds70lWePNU7Ect4QGJppZlnmcaKI6wG7sHQVGaKDavyvR8tzvR6K3ksgUotnLOun1eBAPZ
OoD25wI6vescDnyA7zKuVoDIjnuGqg6QwWNwaFUH9tQ2CGXlgnApuoxNxtF7dPMXNpBJeknXuSP1
akXsJvsUEcG4TZwxorlxI6jV3+3/5pxUdQ+6Vj1+ufK970kQhUguKl3TNxJorTZkTtHLom3W3rAU
jJvuZgVlauCz6w8vnqc0IFkhQj0BnU4LVp3LFkrZpiq9YP4C1JsQ8XQk3H/gEosPYeelBvlP0Fr4
Czlm0DJGWGFuC/NtTdomHo1UC2pkYoWHSPactB8y2hRYhufqJC1cYLqgaPAJi4C+dCGMFpjyTLyy
ysF7LzSMVGanS7DpLE1r6TPgalbu/G12Ozsj7s1nB/ElgKorkTkhi4Df7nDwUD7Kv7CCy4pcO9as
BKKMs8czPPyWbFVl6DkMBICYkfXnwsALTpi2c4jAZ5wOgC9V3STDlk4Q34RwM6o/YGss831X3TkZ
EiXew3j4OnAt4xk8Lp+u6c2lH/MFlcXqp4XMjcMCTBYr+NoZ2YNO5h6ObCT7YEWzQw8wY81SDZ1m
knA658CPKBosP0MYwcDajMsiUrXEUS1oeRN0OghSk78ixXFpLuI5OHRzDrLTnreCXD59+e5wOkTF
a1E4GYak9uk0fPARiVi3ksXe2/SsBc5fAJHhSKmsQDcLchTzQqxh/Wof8mkwQVw/1SdxB1KMjNod
3oo7DOqgucNcolYrelHBGb058ibGl1G9ZbOr3o1sTrkeSRCBlrDSzRScCcm2O2LgtxnoB+U15O/a
4KP23m2qGkvBt5d/CngShsJi/KLnhSostPWaAO59I7zsKAoDjlNi3XhVLqKicj0qzUvG4FyfF6Uw
2YdomkvktZyv4fcEwsGkle+Cfj/71nL9wCbbErqisKfA5SPIpxnDo0PBrjZiKpA9eD9o57/ANyov
OhKoSpnilI/XVtYLAVkiC+z3YUb0Syp56Kg0n5Qqr3MATykZjmIckrdQ7Wvk6RnA87qZrAVb+VAZ
iqew/mRKxUr7AUTzHT++DLfyMv3bLePnZ+ia6YcxMh+UagVXsvKCCSUeMuCerp/tP6ZQJGmDnNWs
/IsokGhNRnWOJ2O7pVHQ4+nP3IcvBLk2WcUn2n4GJCMk728POElieFecag1n1aqiZ2pX9CU3o15e
T0cCgvZw2xMmgktqpRGtlnlpl6pMx2x3p6Yx5tTQsx7Zem2zJkVs3P2QtYu8+sz4eSnKXgNLZQwG
qFImu0M3Lhe1eZ/eBG440fpjoOzE3thgmsXbzh4f/zEh7RRq9zb/1PRW+FVJaziqXYhfIRXZaNV9
ZvXHklPrmleYNXT+Bf/ZuWJTOG3HEQvArVE0CKwwm9bSmHrGGqBVjarjfunemJSuxs29XUPgQ1BY
tvgIiDoYSntq/QIBRh48C2HzG96iM65GxmS1oiO3/Qlk83OgN88RMvmJT+iwAZwianVwz8WstNhU
QcusSkal0P5zvaxb34x/32yBaKSX08ABQdBNyngcibq+Wt3tRT4YTYieWa0Wh8s87oEMjIibep0p
KS4qocQ/T7KYP16uPkF4S1hFKpqefJmAuSBvBgJVYTodgND2OUoLLbtTzl9V/mhcDyl8jBbWwdPm
6bwxQ77nAb1eK627RKSuFuTnEjlrU71M45hEri+qZL5D5wZgsCqh+TUvedp7acQqH3H3yD+tRYRg
xxpY6i9BQFubdryF3V+t19gpS89NmCNVNgCszMHKlV7crownKJGGzAKipg9cs8TVm0IfYzU4mkRB
iUQhvqpNl3cPZHAbnfHed0gaYc6Zn4PfUwQv5BPAcNfQZURwuT69sJ2A9Wp+sjMDh5EDlN7j71Rq
rOTPqkCTIrXhrNxatHOJGYhr+suCAQk0oMZz1jlzruRw1o/NvrBFSFlQSaRUqmTr7yJQ4sgv6RA6
XbGMfip6O672lGcYt11faTC+wIjf2YDtDkFGDirdGJ3r+X4+JX3PwOkLdR9eKjTysniDnb8L26l7
vnMYYTbSHTA4hAtGnatogLRWjTPVwzEH31DBwZiElNjTPmFy8BIIbeK+kII+dlK5L5+rKywPv/yc
ROYp7OevCHgy5vU/17RCWi5nEc35HDmJDUKXN/tM6S97qr+hOaE8ToljVP/EESjGgvygVRZaH2Bh
jQHL8DxoHQzDZvlu5k3mfH5GseJvSEbk6PiM7wNJ8AEbYfHTIRLVgf/Ifk69FlrGm6m87VeiVOTI
5KKkeE90nkVssSgMrTilLmN1vB82VTmFseOyKaDk5FY7D4GZjMHM6adc6CXgqmoIaOPGW5i1957i
8qMh/WsZpgLh8t7vo/+aO3cwjGGxw2dPy8TnqNwfBxSAKWf1/F4nLJBslWcHiry4P0cVcnac9ETI
68XCAUYezfUcTlTQjJGOpZNeiMPAErkzv9DfWHRSxcIvv8pcUeLWUsnC8WSY0Oal47h4HSbpIlrZ
R0hHfN21XrOCulP/Jvi1KvVho1PLoX6pb9yWTAthBOp4uNFr0lJXX5WuZXqvfPnB0CRWyW21x3ml
qkOaVYrDui46UCCMI8o19v00esYdPckNlcorrcZuJVnYb0WgVqFlllRrlRv93n6muoDKXi1hrAxt
rtaAO8VtC3wwz6NWtG5ibfGywDsOLM8vs9DH859jrBZ4R7jYdtucdWjkWV5E3i8Ria6c9qp4ROeL
jfSvpfleBzb3bkwI/alMmdvjOlYfWUJoRrcTSkZlOVGpXxaUkhObKpr6ZuIqhdaR1kk6YmlqtAMx
LfWSQEL9Ywo8yxx9yC16lj9AeBnfojOD33cirhWNRDi1ErNM8VuvqNuToBnRqv2gSZ1o9Sxz9kB7
p5peK7UwszBHA9pySqLnd6bsATpKeJKjj7FtyBt0ynHlUicqOMtThhZlSc07z/d3EzdOtN9ydC7B
jG8dOwV9UaVUHPdTiw+/yZ25TIA/JDZAOFr9oLpsNW8+5dPZynaGZ2nBv0vsxTaq0WPNgHxUiS0c
8LaWFLtwRKZOr6zN9l8JzIGMsAspk4Rk1aL8XernDlU2AAdqqmm+Qd4MWY4xw88f73ZwOswOK4Lz
9mu4WDzMB9rhs9zHLVuHKNZsGDoC5ntHpF03AeFveNopGaxfGVmJUZmMVjYIQsH3aEvz3LiUI1Hu
MUevM8LtvBjikGWZ2VBWCYS7YBGDHRao7TOYF2gltNp5rhKLTtEuZ+tstJYKRb8qpipv0djidJbf
A90BdQltGeymKVkZ97dDLEmi5gbPeMgWuIZL0J4Ee3YNA2cctXPJ+v+NRtTWa70Qvzy/lxobOs6D
abonwLpm1BgKnNySbeRvYgIdj3X8sT85ht2CqJv+xmozAXcpOInOTPzbW8jQTjkOWXkd2z6svnkK
b7r+d53LJSH1puNR+FGr0tZymWfZ1qnVBW/svUYRAoEDwEZpu0gxFJpS4znf0aYheSZ7LRQqVWz9
t9ZG+WgBAx3n2XTDVM8527ptsloMIL1jrNbWpn0juvKhU+eaYKSs1opH6B8ZCaN8r2fEqoOmNXFN
wqFZuQIBGLnX4AbORvpBhOeDxzzXNau6hZa3NbvcRCQ/IFiPF3J/htnFB9cF2hOtdEJoIGL3PPIs
retoeSIVfXswb8xL3soap9fLMq+f6BuN8t6xDW44104cKMYh8n1bHXWBZEX114rqYPPNVnyiBge9
JlqYVNlEp/IGgBCGrbgYRCPngQwZDphtlDILIkxF0hLOAhVXKlU631B8Q8zTy/ksUNNWJNQpVujA
lLXCT+q7AwSHSTRn+9r5Gw8W3G6a1lBwEtWKukektY8M/1W4TCkao8b1j79br//vFMg9IZTptVev
SpACrTErme50pMl/Xrhie41y7jh583pBNHCyqsICC+2NlyZMcSpaCXevQIc040+hW22lF1N+d3tF
neOm1TzpDILWXUEoINSUexWP/6dIvV/SkInAlVlGXySQ0qOnTHRQlwt5oPaC+pQBXA4J8YMCAKZi
O5HDyw2YrqcYfZYuvuSbJvGrTcGZOwR1bYRPm8h0ye/RnPxvmhYfQjzGktLMcGP1lEIIQfGcCIeY
0h8QrJ7bdsPpEHAzmVRlpPLmra2Cf1BGdcXH4+Wpo62OFCHv2H3Jo/wSJlYMCZaR3ROThUvsqyiU
AEkVugCuuN1UWNuWwy5TvY+qmQ5e/RCcx4hF/S2LzC4rIk86jYGJ+Jb/GTilBenyu/zSovM2xi8a
0oc4Bm+kP2532Jy3l72EdhOqW1evQyNX0+49uxTqqUhjI3XMFvTnd0N+RGXrbEvHD6ueOrML2hoK
Pn6T4BWPFHle1FzN0h2MWlA3LMuaePIs977VtqnCuzx41se/CgcBs9rKwXleJg+ErYhKEv0nvVtc
tgedL+5zsH+GLxC1V8v/qP3GS29aWpZNUZLTcOiFzalwbqkO14kMC4Xy8aPBm06u5feJv0SyOOcN
5tXAYKWlMN5DlAZeJuMVdegRd/IDoiZzGT7HIWj5aAk9oOeCobQs7pswcMcwAtJ1tcAHn2pLYbEW
ADEZpeFJ97j3hSc7boKVusnt6HBsedZBmePcnHjqZwmst8YPb3N8VZOZjId9OpQgapOVDOFyf0SU
DSiv3WM8BSYqlFNTolngBVdUGyEq5Ukg2U8nj2byH0Hax71sbMDfJY1LTqM8HN7wjHkBkwpwBLrQ
a5C+E6+TRbCRUvneKG9OigGAnWvzBhrG3Wigze7vD2QWVGvT6VL+h1XJVuEmGu0Vg/qA0wSxjQv9
QWM9VVMW8aJV37yhiN/JP3dzM1kqFXiGqTNmpBKpc6AAcMm3KmR/RpQk8x5vgu9R1mdK/bXhsK0+
MckJcAJEMhTo6SZODbgT+CbnUNbUCFxTawvGvK0Kgqm2XizqUUSXmcixGgHOK8msH2ptb6jSF6QJ
jKS1wfOC7j0RvCzyLelKFW9JOwYDbkSUR+eMceyiVZpPj4U7Y6PZB0Ov3B6Hgc6TTImsiCC9TIuc
lOavl3HMEeeT6gJko5M5sk48r7Fyp3OCUudcClDNWzq+yzdFsKkBQxPgoibeNWtoWwW7SSvts5lF
Nvrs3LidGwZXf9YNuLDbLCr08jXg4zGFHCo1VjlBrtuh6BJv18tgdqeYaDUhnNFfruvzDcCHbgJr
UdlmLWZ8sEHG4cvWp8Kf0xhJH/kSN5i7PCBchcld5/lpqraObC/TK7llmLkop9OJaxpJcNzVN0H6
87CuUN2YmOQbPy7KECorBsERpGOBQ7w15Vfg839n55tG/wB6yYnGSr50KUEH/5UxgrcrhxQahIHy
DGG1fNymWMJToQdobN/9jvGaGJmUSys/TDyPWnjA8pDS0zXW3YKT5EQhcwh4qpNb56Z4u7lNNJ48
oaj75MNSnXSXczthoaqZIbQ937UUlNTNoinfxeD4rP6hzacFUStW+oIttv3BVg7BFgMH1if09jgz
Eh/ZZ7evEtKbeP4/unM6iDNzCVTJN6shWfiaTeuY991gt9WqaSbTKI+fdwhMCroBXDpwIu7D8cnc
AzRPEfxgN+M8voi9e9RTziULDvENeUSyAKBUAltAWhWFqwa+xyMb2ChxKDJ2pSf9O6uS1yN0kmtp
2dJeM/zdk3zD1p3k2UJV/soJLrbWvDCNQRL0l+OVPLZRJhp2c2Cj5YcsaKO+NNf0TPhXctg4BcLh
nKAS34OaZZTu2evZwqTc+D/qnJgc2COlsmYuHV/YQZzpPM+6KQ8hGNJu+iHBBbEkRc4GnfOYzJda
X3cEoP2KVzloJYG/J25GHqU+kd3gbgaF1SzF0i5MWkzbJ0NWWEXWuLmLuLoOwsFMj4tbPAw07M+4
Ee8R4F47ml13RTBEp8ZiT6LV98tzTjcbcg1QQG8voZ4AP+xw5E59vh3UNXAcWo7YG+ISTNwP9du7
x447UIUatucA3ylV12zum5e33CwZezoiVOq4hornfPSlJIcd6vC4I84PLjp5fOpLL8VIO8OEDTEJ
Q736lPoqslqDPmDPiRQbt6N2ya8zYtMvOUKLWNMrw70JcP5xh4y8/tkdPzZW1PczUmuy4KjG+C/b
ImXk5qsncgDQb4UGKCUWk3v2jUWM4I3GZOxiw8EH7dRdqC/3O2WeQJK+ne7IPvi30XWvSpJx2mv7
AOyWuw/9d990Mi3HDMNmlPzH9GRcYl4afXWNoxN7UsIplBEVr8klOA0CkDq+oUGLQNwp1shakO7l
40eNfpYSKVzOEEWLS6IKxvALTFYP3D0rkxHMCrj+OLUWb+2uRI9bynYarsHdREocYte93gCv5A/T
MBddwUAInDZJzntZWB5r9fmF+z4yZEK/PKd9Ym8vCpBlvy4LHP1hRo/mEo3Odp1FkWZfgBj+0KKh
zXCH7Sa9aq990dIL2ccqwuN+NsWW1wc+1hA8i+pIuYh7KQkzloYklATLYxD92QHOSFUuTL+27u/l
Yj0BZZb4Nu2+BuMtmjeTapMI5C8NicJfVTjCGcfV8iuuhMt+TK2lj7Sm1m32hZdVSCwj0KN81+XI
iOjF3uI/5yU0fr0pnHP2PpPnJ6CkuB724T0nxMOOUG4jM8twrXI7xEKWPhwGMXkzqatGTFzz7vD6
IMouBOBW8bZV6UYo2Za3Ht508NAk8l1Cu5pcfzUixXlruhcd8Hn/pWNPLFx33HxjpOlZbqNf0ZKz
L4vpTMGBzW/kcafBD54nVtNN0Z9Ju1+NAqmW3YbvR1KTt6UHohYefQwXg3sw9W1FK2Xv20U3Zr6D
Igsjik1OKGo77y7hJBCf+3kOFCVsBby+MOnvLK7P6ynNvpy0wqnWCbu+Rn3Jv36eYOCvRftdOJl4
0HNf8pmKlvEz37QNS8fM46kWB4rStBTw5rNeYhpiAn9q/Kb3UTEdNmvm4ecaxECbkAm531n/Vt+l
6cJBdUOoFRWMKWwsBS0Ggsn2lksgauwHjCj76TDFx6L/utCy2ihNYkyYtfdG8dkqPsTe/oPN+OO8
m98jKA0buB8dBVFvI7XJ0POkubNEH33ibM79gS00Agqep064utHLYtbrebeeIAuevk3huCSJPGcO
BBxnCSqBAmZCpparI9+mUtgi1s5NBNrzw8sIeuU/D+TLqBKCxeGWFGB+QI9ZZcpRKeTMmuRh5Hhr
ri+Y4Viz2l0OPZd7wxAFQVqvfXCa3AQlaYpHeh71OLS+bGGrI0WItUk0PtXgzDt9x4WXqV4cROo/
12nFdquGr3OvQEX0+RyeCkTPq/gWXXIsBk0yLQrKJ9zjwzGQJ2j1QYAXDummbHsotrxNtpUUBTpp
PscGuplXfldkScGalsXGrwjLnlZ/RCrqW02xPw0/niB5umCHnQKl3pWKB65XOcUk3/Vln8y0EPpR
e88DEIsn+wk+Fuo0POAvD+CAWns8qKv7kG6cyb5K1Xdl7FAkrzUqTfI0yDsEHGbnDsQRw0+1Rrb+
MYCmtnxBmRbu+GUjQ1BIpUtYJRf5jUOJ7jW9Z07c0oD69h3Qmazo5QrGLowYlGV133Zw1Ccah/Jq
F+IfOsPcw4J8LoKAhYkA3GbASC7qTVy0jGzYksBhJfOSUN0EX2F/m4Vy8UjYTEkV6VYBlgLXVyBY
Qtqj77FSiBNoi5Dm+QSCFarnEelA/wBiFwZcqcSqlmIF62weL358Zy15Otmt94ZOsGhv8siGydSv
QXdOxkn3jfo1Vx3XmhPponJLpfoRaIWyV5dVS1LL/zuF/Xk4ry2clKvdGi8QP8sIAHRhk5GmG+1g
liE0ZBNKZgmVWotp6Ho6tFAV0qcu38+I6UwOEzKEJII4wrgcCc5gr7x54m1/vmuTdWdoWJFlKHqR
XsGGahUd83D8chYeFexCQjUI1V4kce+yrz0WRjFrRYOX6zt+azk3bo40ac5BvqDBlaK6PQbu/Vtb
OoP/J6Pe5S+PJJMFAbjNjvb80FBzeF0oPhu/RwpNodYp01e64JqSMutrTmsFpbJ46t8GsRp4KRqE
Lp7lsxMr4OarWQx25KF8xwFr5ihs99PDiNSaxRT2EPfjYze9NK9fN9mZfW+LuTWwUQOz0fGIerXM
veHwN21w/B18aqXezzSxCKr01XbCdW6VMmd6VvKA8mLqfe3nbFDs0FdIOK0Y9Z/5AbrBRUokGgTZ
gJp1+LRiNnk35U1eKcnZOD3yVqNE1/fYwr1B5/SDiQlXsI8al37fa7gFeTAvoksSQBh2jXAksErD
je1sSwOLkTyQOR0zlcw1O3C55jPGO7n+sJUsrPSTqMTfS0TirvXJs+Y35mqQr0hOfvJkxg2XSulU
OJ05BVZbrG6hHAGqsQUseou632u7870ejv8glL9WYbUMQLj4fDRjHkANEXjD6SIoXjtgtxk29yl3
X9cj1D3jxHJeaNXlXET6FUfkHYd+JKhAOt9py9MSo4OnykuDbioBWFBHdut0V253SRhrpizuFUne
5O3JXSTSYvLhFHg94byt2EcZJN1awBOJ1bQedQcbe7cUokK6QPFwnM54liJmbXhKPxhbc+//MaD/
2eB8GPvC3rzrq1e7
`protect end_protected
